-- code generated from the following source code:
--   ../vm/fail.ecl
--   ../vm/value.ecl
--   ../vm/ram.ecl
--   ../vm/frames.ecl
--   ../vm/vm.ecl
--   ../vm/main.ecl
--
-- with the following command:
--
--    ./eclat -arg=true -relax -notyB ../vm/fail.ecl ../vm/value.ecl ../vm/ram.ecl ../vm/frames.ecl ../vm/vm.ecl ../vm/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute1875, \$127_copy_args_to_heap544\, \$128_pow568\, \$129_div569\, \$130_mul570\, \$131_sub571\, \$132_add572\, \$615_forever5741837\, \$640_forever5741836\, \$665_forever5741835\, \$689_forever5741833\, \$698_forever5741834\, pause_getI1880, pause_getI1890, pause_getI1898, pause_getI1906, pause_getI1914, pause_getII1881, pause_getII1891, pause_getII1899, pause_getII1907, pause_getII1915, pause_setI1876, pause_setII1877, q_wait1878, q_wait1882, q_wait1892, q_wait1900, q_wait1908, q_wait1916);
  signal \state\: t_state;
  type t_state_var2552 is (compute2415, \$400_copy_args_to_heap544\, \$401_pow568\, \$402_div569\, \$403_mul570\, \$404_sub571\, \$405_add572\, \$462_forever5741867\, \$466_forever5741861\, \$491_forever5741866\, \$495_forever5741861\, \$520_forever5741865\, \$524_forever5741861\, \$548_forever5741863\, \$552_forever5741861\, \$561_forever5741864\, \$565_forever5741861\, pause_getI2420, pause_getI2430, pause_getI2438, pause_getI2446, pause_getI2454, pause_getII2421, pause_getII2431, pause_getII2439, pause_getII2447, pause_getII2455, pause_setI2416, pause_setI2460, pause_setI2465, pause_setI2470, pause_setI2476, pause_setI2482, pause_setI2487, pause_setI2492, pause_setI2497, pause_setI2503, pause_setI2508, pause_setI2513, pause_setI2520, pause_setI2525, pause_setI2530, pause_setI2535, pause_setI2540, pause_setII2417, pause_setII2461, pause_setII2466, pause_setII2471, pause_setII2477, pause_setII2483, pause_setII2488, pause_setII2493, pause_setII2498, pause_setII2504, pause_setII2509, pause_setII2514, pause_setII2521, pause_setII2526, pause_setII2531, pause_setII2536, pause_setII2541, q_wait2418, q_wait2422, q_wait2432, q_wait2440, q_wait2448, q_wait2456, q_wait2462, q_wait2467, q_wait2472, q_wait2478, q_wait2484, q_wait2489, q_wait2494, q_wait2499, q_wait2505, q_wait2510, q_wait2515, q_wait2522, q_wait2527, q_wait2532, q_wait2537, q_wait2542);
  signal state_var2552: t_state_var2552;
  type t_state_var2551 is (compute2412);
  signal state_var2551: t_state_var2551;
  type t_state_var2550 is (compute2407);
  signal state_var2550: t_state_var2550;
  type t_state_var2549 is (compute1922, \$117_forever5731839\, \$117_forever5731846\, \$117_forever5731847\, \$117_forever5731848\, \$117_forever5731849\, \$120_forever5741838\, \$120_forever5741850\, \$120_forever5741851\, \$120_forever5741852\, \$120_forever5741853\, \$120_forever5741854\, \$120_forever5741855\, \$120_forever5741856\, \$120_forever5741857\, \$120_forever5741858\, \$120_forever5741859\, \$120_forever5741860\, \$143_copy_args_to_heap544\, \$144_pow568\, \$145_div569\, \$146_mul570\, \$147_sub571\, \$148_add572\, \$149_vm_run_code547\, \$208_forever5731845\, \$212_forever5731839\, \$258_forever5741844\, \$262_forever5741838\, \$287_forever5741843\, \$291_forever5741838\, \$316_forever5741842\, \$320_forever5741838\, \$344_forever5741840\, \$348_forever5741838\, \$357_forever5741841\, \$361_forever5741838\, pause_getI1927, pause_getI1937, pause_getI1945, pause_getI1953, pause_getI1961, pause_getI1984, pause_getI1995, pause_getI2006, pause_getI2017, pause_getI2028, pause_getI2039, pause_getI2065, pause_getI2069, pause_getI2094, pause_getI2105, pause_getI2116, pause_getI2123, pause_getI2130, pause_getI2142, pause_getI2149, pause_getI2161, pause_getI2177, pause_getI2188, pause_getI2199, pause_getI2215, pause_getI2226, pause_getI2237, pause_getI2244, pause_getI2260, pause_getI2271, pause_getI2282, pause_getI2290, pause_getI2303, pause_getI2307, pause_getI2314, pause_getI2321, pause_getI2329, pause_getI2337, pause_getI2348, pause_getI2359, pause_getI2367, pause_getI2375, pause_getI2386, pause_getI2397, pause_getII1928, pause_getII1938, pause_getII1946, pause_getII1954, pause_getII1962, pause_getII1985, pause_getII1996, pause_getII2007, pause_getII2018, pause_getII2029, pause_getII2040, pause_getII2066, pause_getII2070, pause_getII2095, pause_getII2106, pause_getII2117, pause_getII2124, pause_getII2131, pause_getII2143, pause_getII2150, pause_getII2162, pause_getII2178, pause_getII2189, pause_getII2200, pause_getII2216, pause_getII2227, pause_getII2238, pause_getII2245, pause_getII2261, pause_getII2272, pause_getII2283, pause_getII2291, pause_getII2304, pause_getII2308, pause_getII2315, pause_getII2322, pause_getII2330, pause_getII2338, pause_getII2349, pause_getII2360, pause_getII2368, pause_getII2376, pause_getII2387, pause_getII2398, pause_setI1923, pause_setI1969, pause_setI1973, pause_setI2044, pause_setI2049, pause_setI2083, pause_setI2135, pause_setI2154, pause_setI2166, pause_setI2204, pause_setI2249, pause_setI2295, pause_setI2299, pause_setI2325, pause_setI2333, pause_setI2363, pause_setI2371, pause_setI2391, pause_setII1924, pause_setII1970, pause_setII1974, pause_setII2045, pause_setII2050, pause_setII2084, pause_setII2136, pause_setII2155, pause_setII2167, pause_setII2205, pause_setII2250, pause_setII2296, pause_setII2300, pause_setII2326, pause_setII2334, pause_setII2364, pause_setII2372, pause_setII2392, q_wait1925, q_wait1929, q_wait1939, q_wait1947, q_wait1955, q_wait1963, q_wait1971, q_wait1975, q_wait1986, q_wait1997, q_wait2008, q_wait2019, q_wait2030, q_wait2041, q_wait2046, q_wait2051, q_wait2067, q_wait2071, q_wait2085, q_wait2096, q_wait2107, q_wait2118, q_wait2125, q_wait2132, q_wait2137, q_wait2144, q_wait2151, q_wait2156, q_wait2163, q_wait2168, q_wait2179, q_wait2190, q_wait2201, q_wait2206, q_wait2217, q_wait2228, q_wait2239, q_wait2246, q_wait2251, q_wait2262, q_wait2273, q_wait2284, q_wait2292, q_wait2297, q_wait2301, q_wait2305, q_wait2309, q_wait2316, q_wait2323, q_wait2327, q_wait2331, q_wait2335, q_wait2339, q_wait2350, q_wait2361, q_wait2365, q_wait2369, q_wait2373, q_wait2377, q_wait2388, q_wait2393, q_wait2399);
  signal state_var2549: t_state_var2549;
  type array_value_68 is array (natural range <>) of value(0 to 67);
  type array_value_72 is array (natural range <>) of value(0 to 71);
  type array_value_128 is array (natural range <>) of value(0 to 127);
  signal arr1868 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1868_value\ : value(0 to 67);
  signal \$arr1868_ptr\ : natural range 0 to 99;
  signal \$arr1868_ptr_write\ : natural range 0 to 99;
  signal \$arr1868_write\ : value(0 to 67);
  signal \$arr1868_write_request\ : std_logic := '0';
  signal arr1869 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1869_value\ : value(0 to 67);
  signal \$arr1869_ptr\ : natural range 0 to 99;
  signal \$arr1869_ptr_write\ : natural range 0 to 99;
  signal \$arr1869_write\ : value(0 to 67);
  signal \$arr1869_write_request\ : std_logic := '0';
  signal arr1870 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1870_value\ : value(0 to 67);
  signal \$arr1870_ptr\ : natural range 0 to 99;
  signal \$arr1870_ptr_write\ : natural range 0 to 99;
  signal \$arr1870_write\ : value(0 to 67);
  signal \$arr1870_write_request\ : std_logic := '0';
  signal arr1871 : array_value_72(0 to 99) := (others => (others => '0'));
  signal \$arr1871_value\ : value(0 to 71);
  signal \$arr1871_ptr\ : natural range 0 to 99;
  signal \$arr1871_ptr_write\ : natural range 0 to 99;
  signal \$arr1871_write\ : value(0 to 71);
  signal \$arr1871_write_request\ : std_logic := '0';
  signal arr1872 : array_value_128(0 to 99) := (others => (others => '0'));
  signal \$arr1872_value\ : value(0 to 127);
  signal \$arr1872_ptr\ : natural range 0 to 99;
  signal \$arr1872_ptr_write\ : natural range 0 to 99;
  signal \$arr1872_write\ : value(0 to 127);
  signal \$arr1872_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1868_write_request\ = '1' then
                    arr1868(\$arr1868_ptr_write\) <= \$arr1868_write\;
                  else
                   \$arr1868_value\ <= arr1868(\$arr1868_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1869_write_request\ = '1' then
                    arr1869(\$arr1869_ptr_write\) <= \$arr1869_write\;
                  else
                   \$arr1869_value\ <= arr1869(\$arr1869_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1870_write_request\ = '1' then
                    arr1870(\$arr1870_ptr_write\) <= \$arr1870_write\;
                  else
                   \$arr1870_value\ <= arr1870(\$arr1870_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1871_write_request\ = '1' then
                    arr1871(\$arr1871_ptr_write\) <= \$arr1871_write\;
                  else
                   \$arr1871_value\ <= arr1871(\$arr1871_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1872_write_request\ = '1' then
                    arr1872(\$arr1872_ptr_write\) <= \$arr1872_write\;
                  else
                   \$arr1872_value\ <= arr1872(\$arr1872_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$397\, \$136\ : value(0 to 1) := (others => '0');
      variable \$403_mul570_arg\, \$127_copy_args_to_heap544_arg\, 
               \$132_add572_arg\, \$129_div569_arg\, \$146_mul570_arg\, 
               \$130_mul570_arg\, \$144_pow568_arg\, \$147_sub571_arg\, 
               \$401_pow568_arg\, \$400_copy_args_to_heap544_arg\, 
               \$404_sub571_arg\, \$402_div569_arg\, 
               \$143_copy_args_to_heap544_arg\, \$148_add572_arg\, 
               \$128_pow568_arg\, \$405_add572_arg\, \$131_sub571_arg\, 
               \$145_div569_arg\ : value(0 to 95) := (others => '0');
      variable \$v2139\, \$v2379\, \$v2120\, \$v1942\, \$v2053\, \$v1903\, 
               \$v1988\, \$v2098\, \$v2451\, \$v2054\, \$v1934\, \$v2443\, 
               \$v2230\, \$v2341\, \$v2352\, \$v1968\, \$v2087\, \$v2219\, 
               \$v2253\, \$v1895\, \$v2181\, \$v2275\, \$v2057\, \$v1178\, 
               \$v2060\, \$v1977\, \$v2435\, \$v2109\, \$v2010\, \$v1999\, 
               \$v2170\, \$v2021\, \$v2427\, \$v1950\, \$v2241\, \$v2264\, 
               \$v2146\, \$v2032\, \$v1887\, \$v2208\, \$v1911\, \$v2192\, 
               \$v2127\, \$v2311\, \$v2158\, \$v1958\, \$v2294\, \$v2074\, 
               \$v2318\ : value(0 to 63) := (others => '0');
      variable \$191_instr\, \$v2395\ : value(0 to 71) := (others => '0');
      variable \$v2381\, \$v2210\, \$v2194\, \$v2221\, \$v2001\, \$v2183\, 
               \$113_p\, \$v2034\, \$v2266\, \$v2232\, \$v2012\, \$v2100\, 
               \$v2089\, \$v2518\, \$v1990\, \$v2172\, \$v2023\, \$v2255\, p, 
               \$v2277\, \$v2354\, \$v2111\, \$v2076\, \$v2343\, \$v1979\, 
               \$v2286\ : value(0 to 4) := (others => '0');
      variable \$v1944\, \$v2278\, \$v2112\, \$v2222\, \$v2077\, \$v2080\, 
               \$v2396\, \$v2187\, \$v2002\, \$v2024\, \$v1905\, \$v2267\, 
               \$v2236\, \$v2184\, \$v1936\, \$v2256\, \$v1913\, \$v2005\, 
               \$v2243\, \$v2233\, \$v2104\, \$v2062\, \$v2437\, \$v2122\, 
               \$v2016\, \$v2445\, \$v1889\, \$v1960\, \$v2355\, \$v1897\, 
               \$v2038\, \$v2093\, \$v2270\, \$v2141\, \$v1980\, \$v2013\, 
               \$v2382\, \$v2101\, \$v2320\, \$v2160\, \$v2211\, \$v2453\, 
               \$v2195\, \$v2027\, \$v2313\, \$v1952\, \$v2148\, \$v2198\, 
               \$v2429\, \$v2344\, \$v2176\, \$v2287\, \$v2225\, \$v2358\, 
               \$v2115\, \$v2056\, \$v2214\, \$v2090\, \$v1994\, \$v2289\, 
               \$v1983\, \$v1991\, \$v2173\, \$v2259\, \$v2347\, \$v2059\, 
               \$v2385\, \$v2035\, \$v2129\, \$v2281\, \$v2064\ : value(0 to 3) := (others => '0');
      variable \$149_vm_run_code547_arg\ : value(0 to 294) := (others => '0');
      variable \$v1701\ : value(0 to 127) := (others => '0');
      variable \$v2501\, \$v2516\, cond, \$v2075\, \$v2031\, \$v2218\, 
               \$v2209\, \$v2545\, \$v2097\, \$v2052\, \$v1918\, \$v2463\, 
               rdy2414, \$v2191\, \$v2252\, \$v2231\, \$v2317\, \$v2268\, 
               \$v1987\, \$v2072\, \$v2543\, \$v2380\, \$v1941\, x, \$v2153\, 
               \$v2400\, \$v2014\, \$v1976\, \$v2157\, \$v1910\, \$v1930\, 
               \$v2310\, \$v2022\, \$98_a1\, \$v2404\, \$v2223\, \$v2362\, 
               \$v2389\, \$v1931\, \$v2276\, \$395\, \$v2324\, \$v2174\, 
               \$v2234\, \$v1885\, \$v1965\, \$v2152\, \$v2336\, \$v2507\, 
               \$v2078\, \$v2086\, \$v1948\, \$v2229\, \$v1972\, \$v2345\, 
               \$v2423\, \$v2332\, \$v2240\, \$v2169\, \$v1932\, b2, 
               \$v2003\, \$v2293\, \$v2196\, \$v2033\, \$115_b\, \$v1957\, 
               \$v2401\, \$v2182\, \$v2479\, \$v2126\, \$v2025\, \$v2425\, 
               \$v2441\, \$v1966\, \$v2119\, \$v2351\, \$v1926\, \$v1902\, 
               \$v2274\, \$v2138\, result2413, \$v1893\, \$v1901\, \$v2485\, 
               \$v2533\, \$v2353\, \$v2108\, \$v1894\, \$v2433\, \$v2442\, 
               \$v2298\, \$v2285\, rdy2406, \$v1919\, \$v2185\, \$v2000\, 
               \$v1964\, \$v1998\, \$v2370\, \$v1989\, \$v2247\, condition, 
               \$v2495\, \$v2500\, \$v2165\, \$v2113\, \$v2047\, \$v1884\, 
               \$v2073\, \$v1879\, \$v2366\, \$v2523\, \$v2394\, \$v2546\, 
               \$v1886\, \$v2374\, \$v2356\, \$v2164\, \$v2202\, \$v2426\, 
               \$v2468\, \$v2011\, result2410, \$v2220\, \$v1940\, \$v2254\, 
               rdy1874, \$v2490\, \$v2517\, \$v2548\, \$v2133\, \$v2248\, 
               \$v2424\, \$v2458\, \$v1883\, \$v2099\, \$v2042\, result1920, 
               \$v2473\, res, \$v1978\, \$v2263\, \$v2036\, \$v2340\, 
               \$v2506\, \$v2257\, \$v2434\, \$v2102\, \$v2020\, \$v2419\, 
               \$v2171\, \$v2306\, \$v2538\, \$v2459\, \$v2528\, \$v2110\, 
               \$v2279\, \$v2180\, result1873, \$v2145\, \$v2081\, \$v1917\, 
               \$v2402\, \$149_vm_run_code547_result\, \$v1992\, \$v2193\, 
               \$v2265\, \$v2328\, \$v1933\, \$v2449\, \$v2068\, \$v2212\, 
               \$v2048\, \$v2342\, \$v2383\, \$v1956\, \$v2409\, \$v2009\, 
               \$134_is_loaded\, \$v2082\, \$v2450\, \$v1981\, \$v2088\, 
               \$v2496\, \$v2390\, \$v2378\, rdy1921, \$v1909\, \$v2457\, 
               \$v1949\, \$v2134\, \$v2207\, rdy2411, \$v2539\, \$v2091\, 
               \$v2511\, \$v2302\ : value(0 to 0) := (others => '0');
      variable \$v2486\, \$v2464\, \$144_pow568_result\, \$v2474\, 
               \$146_mul570_result\, \$631_int_value\, \$v2524\, scd_operand, 
               \$200_i\, debut, \$482_int_value\, \$99_a\, \$v2491\, 
               \$487_a\, \$v2203\, \$135_cy\, \$114_n\, \$283_a\, \$v2512\, 
               \$307_int_value\, \$193_l\, \$453_int_value\, 
               \$606_int_value\, \$197_i\, \$312_a\, \$199_i\, b, 
               \$278_int_value\, \$v2043\, 
               \$143_copy_args_to_heap544_result\, \$661_a\, \$v2534\, 
               \$v2469\, fst_operand, \$511_int_value\, \$335_divisor\, 
               \$148_add572_result\, base, \$458_a\, \$v2480\, \$636_a\, 
               \$147_sub571_result\, result2405, \$353_a\, \$254_a\, 
               \$196_l\, \$v2529\, \$201_i\, \$192_n\, \$694_a\, \$557_a\, 
               \$195_l\, \$539_divisor\, exponent, \$516_a\, resultat, 
               \$680_divisor\, \$656_int_value\, \$198_l\, \$249_int_value\, 
               \$145_div569_result\, \$393\, a, \$611_a\ : value(0 to 31) := (others => '0');
      variable \$165\ : value(0 to 293) := (others => '0');
      variable \$v251\, \$v2037\, \$v177\, \$v2140\, \$v72\, \$v255\, 
               \$v149\, first_value, \$352\, \$v2312\, \$248_v\, \$v2055\, 
               \$v2444\, \$v1896\, \$v2235\, \$655_v\, \$v1967\, \$v81\, 
               \$v1959\, \$v212\, \$v2384\, \$v1888\, \$v2103\, \$v2128\, 
               \$v2026\, \$630_v\, \$v167\, \$v247\, \$v2063\, \$726\, 
               \$v2159\, \$v75\, \$v263\, \$693\, \$v1912\, \$v219\, \value\, 
               \$v174\, \$v70\, \$v78\, \$v2519\, \$v117\, \$v1993\, 
               \$277_v\, \$v139\, v, \$v2502\, \$v2481\, \$v2436\, \$605_v\, 
               \$v91\, \$v244\, \$v2121\, \$v42\, \$v142\, \$v2061\, \$v26\, 
               second_value, \$v2147\, \$452_v\, \$v2175\, \$v184\, \$v2197\, 
               \$v1951\, \$v33\, \$v1935\, \$389\, \$v2224\, \$v2004\, 
               \$v93\, \$v2452\, \$v2475\, \$v2186\, \$v23\, \$v2079\, 
               \$v2280\, \$306_v\, var, \$v2428\, \$v2242\, \$v2319\, \$556\, 
               \$v36\, \$v1904\, \$v39\, \$v2258\, \$v2346\, \$v2213\, 
               \$v2092\, \$v2269\, \$v2288\, \$v209\, \$v2015\, \$v2357\, 
               \$481_v\, \$v2114\, \$204_v\, \$593\, local_value, \$v2058\, 
               \$v1943\, \$510_v\, \$v1982\ : value(0 to 67) := (others => '0');
      variable \$arr1868_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1869_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1870_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1871_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1872_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$145_div569_arg\); default_zero(\$611_a\); 
          default_zero(a); default_zero(\$v2064\); default_zero(\$v1982\); 
          default_zero(\$v2281\); default_zero(\$v2286\); 
          default_zero(\$v2129\); default_zero(\$393\); 
          default_zero(\$v2302\); default_zero(\$v2511\); 
          default_zero(\$510_v\); default_zero(\$v2035\); 
          default_zero(\$v2091\); default_zero(\$145_div569_result\); 
          default_zero(\$v2539\); default_zero(rdy2411); 
          default_zero(\$v1943\); default_zero(\$v1979\); 
          default_zero(\$v2207\); default_zero(\$v2385\); 
          default_zero(\$v2059\); default_zero(\$v2134\); 
          default_zero(\$249_int_value\); default_zero(\$v1949\); 
          default_zero(\$v2457\); default_zero(\$v1909\); 
          default_zero(\$131_sub571_arg\); default_zero(\$v2058\); 
          default_zero(\$v2347\); default_zero(local_value); 
          default_zero(\$198_l\); default_zero(\$593\); 
          default_zero(\$656_int_value\); default_zero(rdy1921); 
          default_zero(\$v2318\); default_zero(\$405_add572_arg\); 
          default_zero(\$v2378\); default_zero(\$204_v\); 
          default_zero(\$v2114\); default_zero(\$v2343\); 
          default_zero(\$v2259\); default_zero(\$v2390\); 
          default_zero(\$v2496\); default_zero(\$v2173\); 
          default_zero(\$481_v\); default_zero(\$v2357\); 
          default_zero(\$v2088\); default_zero(\$v2015\); 
          default_zero(\$v2076\); default_zero(\$v1991\); 
          default_zero(\$v1981\); default_zero(\$v209\); 
          default_zero(\$v2288\); default_zero(\$v1983\); 
          default_zero(\$v2289\); default_zero(\$v1994\); 
          default_zero(\$680_divisor\); default_zero(\$v2090\); 
          default_zero(resultat); default_zero(\$v2214\); 
          default_zero(\$v2269\); default_zero(\$v2450\); 
          default_zero(\$v2082\); default_zero(\$v2111\); 
          default_zero(\$516_a\); default_zero(\$v2092\); 
          default_zero(\$134_is_loaded\); default_zero(\$v2213\); 
          default_zero(\$v2074\); default_zero(\$v2354\); 
          default_zero(\$v2056\); default_zero(\$v2115\); 
          default_zero(\$v2009\); default_zero(\$v2277\); 
          default_zero(exponent); default_zero(\$v2358\); 
          default_zero(\$v2346\); default_zero(\$v2258\); 
          default_zero(\$v2409\); default_zero(\$v2225\); default_zero(p); 
          default_zero(\$v1956\); default_zero(\$v2255\); 
          default_zero(\$v2383\); default_zero(\$v39\); 
          default_zero(\$v2287\); default_zero(\$v2176\); 
          default_zero(\$v2344\); default_zero(\$v1904\); 
          default_zero(\$v2342\); default_zero(\$v36\); 
          default_zero(\$v2429\); default_zero(\$v2198\); 
          default_zero(\$v2048\); default_zero(\$v2148\); 
          default_zero(\$v2212\); default_zero(\$v2068\); 
          default_zero(\$v2449\); default_zero(\$556\); 
          default_zero(\$v1933\); default_zero(\$v2328\); 
          default_zero(\$v2265\); default_zero(\$539_divisor\); 
          default_zero(\$v2193\); default_zero(\$v1992\); 
          default_zero(\$v1952\); default_zero(\$195_l\); 
          default_zero(\$v2313\); default_zero(\$149_vm_run_code547_result\); 
          default_zero(\$v2402\); default_zero(\$557_a\); 
          default_zero(\$v1917\); default_zero(\$v2319\); 
          default_zero(\$694_a\); default_zero(\$v2081\); 
          default_zero(\$v2145\); default_zero(result1873); 
          default_zero(\$v2180\); default_zero(\$128_pow568_arg\); 
          default_zero(\$v2279\); default_zero(\$v2027\); 
          default_zero(\$v2242\); default_zero(\$192_n\); 
          default_zero(\$v2110\); default_zero(\$v2528\); 
          default_zero(\$v2023\); default_zero(\$v2294\); 
          default_zero(\$v2459\); default_zero(\$v2195\); 
          default_zero(\$v2428\); default_zero(\$v1958\); 
          default_zero(\$v2538\); default_zero(\$201_i\); 
          default_zero(\$v2306\); default_zero(\$v2171\); 
          default_zero(\$v2419\); default_zero(var); default_zero(\$v2158\); 
          default_zero(\$v2020\); default_zero(\$v2529\); 
          default_zero(\$v2102\); default_zero(\$v2434\); 
          default_zero(\$196_l\); default_zero(\$v2453\); 
          default_zero(\$v2257\); default_zero(\$254_a\); 
          default_zero(\$v2395\); default_zero(\$v2172\); 
          default_zero(\$v1990\); default_zero(\$v2506\); 
          default_zero(\$353_a\); default_zero(\$191_instr\); 
          default_zero(\$306_v\); default_zero(\$v2340\); 
          default_zero(\$v2036\); default_zero(\$v2280\); 
          default_zero(\$v2263\); default_zero(\$v2211\); 
          default_zero(\$v2311\); default_zero(\$v2127\); 
          default_zero(\$v2079\); default_zero(\$v1978\); default_zero(res); 
          default_zero(\$148_add572_arg\); 
          default_zero(\$149_vm_run_code547_arg\); default_zero(\$v23\); 
          default_zero(\$v2473\); default_zero(result1920); 
          default_zero(result2405); default_zero(\$v2042\); 
          default_zero(\$147_sub571_result\); default_zero(\$v2186\); 
          default_zero(\$v2518\); default_zero(\$v2475\); 
          default_zero(\$v2452\); default_zero(\$636_a\); 
          default_zero(\$v2099\); default_zero(\$v1883\); 
          default_zero(\$v93\); default_zero(\$v2192\); 
          default_zero(\$v2089\); default_zero(\$v2458\); 
          default_zero(\$v2424\); 
          default_zero(\$143_copy_args_to_heap544_arg\); 
          default_zero(\$v2248\); default_zero(\$v2004\); 
          default_zero(\$v2224\); default_zero(\$v2133\); 
          default_zero(\$389\); default_zero(\$v1935\); default_zero(\$v33\); 
          default_zero(\$v2548\); default_zero(\$v1911\); 
          default_zero(\$v2160\); default_zero(\$v2480\); 
          default_zero(\$v1951\); default_zero(\$v2517\); 
          default_zero(\$v2490\); default_zero(\$v2320\); 
          default_zero(rdy1874); default_zero(\$v2254\); 
          default_zero(\$v2197\); default_zero(\$v2101\); 
          default_zero(\$v1940\); default_zero(\$v2220\); 
          default_zero(\$v184\); default_zero(\$458_a\); 
          default_zero(\$136\); default_zero(\$v2382\); 
          default_zero(\$v2175\); default_zero(result2410); 
          default_zero(\$v2100\); default_zero(\$v2011\); 
          default_zero(\$165\); default_zero(\$v2013\); 
          default_zero(\$v2468\); default_zero(\$v2426\); default_zero(base); 
          default_zero(\$148_add572_result\); default_zero(\$v2202\); 
          default_zero(\$v2164\); default_zero(\$335_divisor\); 
          default_zero(\$v2356\); default_zero(\$v2374\); 
          default_zero(\$452_v\); default_zero(\$v1886\); 
          default_zero(\$v2546\); default_zero(\$v2147\); 
          default_zero(second_value); default_zero(\$v2208\); 
          default_zero(\$v2394\); default_zero(\$v2523\); 
          default_zero(\$v2366\); default_zero(\$v2012\); 
          default_zero(\$v1879\); default_zero(\$v26\); 
          default_zero(\$v1887\); default_zero(\$v2073\); 
          default_zero(\$511_int_value\); default_zero(\$v1884\); 
          default_zero(\$v2047\); default_zero(\$v1980\); 
          default_zero(\$v2113\); default_zero(\$v2141\); 
          default_zero(\$v2061\); default_zero(\$v2270\); 
          default_zero(\$v2165\); default_zero(\$v2500\); 
          default_zero(\$v2495\); default_zero(condition); 
          default_zero(fst_operand); default_zero(\$v2093\); 
          default_zero(\$v142\); default_zero(\$v2038\); 
          default_zero(\$v2247\); default_zero(\$v1989\); 
          default_zero(\$v42\); default_zero(\$v2121\); 
          default_zero(\$v2370\); default_zero(\$v1998\); 
          default_zero(\$v1964\); default_zero(\$v2000\); 
          default_zero(\$v244\); default_zero(\$v2185\); 
          default_zero(\$v91\); default_zero(\$v1919\); 
          default_zero(\$v1897\); default_zero(\$v2355\); 
          default_zero(\$402_div569_arg\); default_zero(\$v2469\); 
          default_zero(\$v2032\); default_zero(rdy2406); 
          default_zero(\$v2146\); default_zero(\$v1960\); 
          default_zero(\$v2285\); default_zero(\$v2534\); 
          default_zero(\$404_sub571_arg\); default_zero(\$605_v\); 
          default_zero(\$v2298\); default_zero(\$661_a\); 
          default_zero(\$143_copy_args_to_heap544_result\); 
          default_zero(\$v2442\); 
          default_zero(\$400_copy_args_to_heap544_arg\); 
          default_zero(\$v2433\); default_zero(\$v1894\); 
          default_zero(\$v2436\); default_zero(\$v2108\); 
          default_zero(\$v2481\); default_zero(\$v2043\); 
          default_zero(\$v2502\); default_zero(\$v1889\); 
          default_zero(\$v2353\); default_zero(v); default_zero(\$v2264\); 
          default_zero(\$v2533\); default_zero(\$v2241\); 
          default_zero(\$278_int_value\); default_zero(\$v1950\); 
          default_zero(\$v2485\); default_zero(\$401_pow568_arg\); 
          default_zero(\$v139\); default_zero(\$397\); default_zero(b); 
          default_zero(\$v1901\); default_zero(\$v2445\); 
          default_zero(\$v2427\); default_zero(\$199_i\); 
          default_zero(\$v2021\); default_zero(\$v2170\); 
          default_zero(\$v1999\); default_zero(\$v2010\); 
          default_zero(\$v1893\); default_zero(\$v2109\); 
          default_zero(\$v2435\); default_zero(\$v2232\); 
          default_zero(\$v2016\); default_zero(\$312_a\); 
          default_zero(\$197_i\); default_zero(\$v2266\); 
          default_zero(\$277_v\); default_zero(result2413); 
          default_zero(\$v2122\); default_zero(\$v1977\); 
          default_zero(\$v2060\); default_zero(\$v1993\); 
          default_zero(\$v117\); default_zero(\$147_sub571_arg\); 
          default_zero(\$v2519\); default_zero(\$606_int_value\); 
          default_zero(\$v2138\); default_zero(\$v1178\); 
          default_zero(\$v2437\); default_zero(\$v2274\); 
          default_zero(\$v78\); default_zero(\$v1902\); 
          default_zero(\$v1926\); default_zero(\$v2351\); 
          default_zero(\$v2119\); default_zero(\$v1701\); 
          default_zero(\$v1966\); default_zero(\$453_int_value\); 
          default_zero(\$v2441\); default_zero(\$v2425\); 
          default_zero(\$v2057\); default_zero(\$v70\); 
          default_zero(\$v2275\); default_zero(\$v2034\); 
          default_zero(\$v174\); default_zero(\$v2025\); 
          default_zero(\$v2181\); default_zero(\$v2126\); 
          default_zero(\$144_pow568_arg\); default_zero(\$193_l\); 
          default_zero(\$v2062\); default_zero(\$v2479\); 
          default_zero(\value\); default_zero(\$v2104\); 
          default_zero(\$v2182\); default_zero(\$v2401\); 
          default_zero(\$v1895\); default_zero(\$v2253\); 
          default_zero(\$v1957\); default_zero(\$115_b\); 
          default_zero(\$307_int_value\); default_zero(\$v2233\); 
          default_zero(\$v2219\); default_zero(\$v219\); 
          default_zero(\$v2243\); default_zero(\$v2033\); 
          default_zero(\$v2005\); default_zero(\$v2196\); 
          default_zero(\$v2293\); default_zero(\$v1912\); 
          default_zero(\$v2003\); default_zero(\$113_p\); 
          default_zero(\$130_mul570_arg\); default_zero(\$v2183\); 
          default_zero(\$693\); default_zero(\$v1913\); 
          default_zero(\$v263\); default_zero(\$v75\); default_zero(b2); 
          default_zero(\$v1932\); default_zero(\$v2169\); 
          default_zero(\$v2240\); default_zero(\$v2512\); 
          default_zero(\$v2256\); default_zero(\$v1936\); 
          default_zero(\$v2332\); default_zero(\$v2159\); 
          default_zero(\$v2001\); default_zero(\$v2423\); 
          default_zero(\$726\); default_zero(\$283_a\); 
          default_zero(\$v2345\); default_zero(\$v2087\); 
          default_zero(\$146_mul570_arg\); default_zero(\$v1972\); 
          default_zero(\$129_div569_arg\); default_zero(\$v1968\); 
          default_zero(\$v2063\); default_zero(\$132_add572_arg\); 
          default_zero(\$127_copy_args_to_heap544_arg\); 
          default_zero(\$v2352\); default_zero(\$v2229\); 
          default_zero(\$v1948\); default_zero(\$v247\); 
          default_zero(\$v167\); default_zero(\$v2184\); 
          default_zero(\$630_v\); default_zero(\$v2086\); 
          default_zero(\$v2078\); default_zero(\$v2221\); 
          default_zero(\$v2507\); default_zero(\$v2236\); 
          default_zero(\$114_n\); default_zero(\$135_cy\); 
          default_zero(\$v2336\); default_zero(\$v2341\); 
          default_zero(\$v2152\); default_zero(\$v2267\); 
          default_zero(\$v2026\); default_zero(\$v2203\); 
          default_zero(\$v1965\); default_zero(\$v1885\); 
          default_zero(\$v2230\); default_zero(\$v2234\); 
          default_zero(\$v2174\); default_zero(\$487_a\); 
          default_zero(\$v2324\); default_zero(\$395\); 
          default_zero(\$v2194\); default_zero(\$v2276\); 
          default_zero(\$v1905\); default_zero(\$v2128\); 
          default_zero(\$v2103\); default_zero(\$v1931\); 
          default_zero(\$v2389\); default_zero(\$v2362\); 
          default_zero(\$v1888\); default_zero(\$v2223\); 
          default_zero(\$v2491\); default_zero(\$v2404\); 
          default_zero(\$v2384\); default_zero(\$98_a1\); 
          default_zero(\$v2022\); default_zero(\$v2310\); 
          default_zero(\$v1930\); default_zero(\$v212\); 
          default_zero(\$v1910\); default_zero(\$v2157\); 
          default_zero(\$v1959\); default_zero(\$v81\); 
          default_zero(\$v1967\); default_zero(\$v2024\); 
          default_zero(\$v2002\); default_zero(\$v1976\); 
          default_zero(\$655_v\); default_zero(\$v2443\); 
          default_zero(\$99_a\); default_zero(\$v1934\); 
          default_zero(\$v2014\); default_zero(\$v2235\); 
          default_zero(\$v2054\); default_zero(\$v2400\); 
          default_zero(\$v1896\); default_zero(\$v2451\); 
          default_zero(\$482_int_value\); default_zero(\$v2153\); 
          default_zero(\$v2444\); default_zero(\$v2055\); 
          default_zero(\$v2098\); default_zero(x); default_zero(\$v1988\); 
          default_zero(\$248_v\); default_zero(\$v1903\); 
          default_zero(\$v2053\); default_zero(debut); 
          default_zero(\$v2187\); default_zero(\$v2312\); 
          default_zero(\$v1941\); default_zero(\$352\); 
          default_zero(\$v2380\); default_zero(\$v2543\); 
          default_zero(first_value); default_zero(\$403_mul570_arg\); 
          default_zero(\$200_i\); default_zero(\$v2072\); 
          default_zero(\$v1987\); default_zero(\$v2268\); 
          default_zero(\$v2317\); default_zero(scd_operand); 
          default_zero(\$v2231\); default_zero(\$v2396\); 
          default_zero(\$v2252\); default_zero(\$v2524\); 
          default_zero(\$631_int_value\); default_zero(\$v2191\); 
          default_zero(\$v1942\); default_zero(rdy2414); 
          default_zero(\$v149\); default_zero(\$v2463\); 
          default_zero(\$v2120\); default_zero(\$v2080\); 
          default_zero(\$v1918\); default_zero(\$v2052\); 
          default_zero(\$v255\); default_zero(\$146_mul570_result\); 
          default_zero(\$v2097\); default_zero(\$v2545\); 
          default_zero(\$v2077\); default_zero(\$v2222\); 
          default_zero(\$v2112\); default_zero(\$v2209\); 
          default_zero(\$v2474\); default_zero(\$v2218\); 
          default_zero(\$144_pow568_result\); default_zero(\$v2031\); 
          default_zero(\$v2278\); default_zero(\$v2210\); 
          default_zero(\$v1944\); default_zero(\$v2075\); 
          default_zero(\$v72\); default_zero(\$v2464\); 
          default_zero(\$v2140\); default_zero(\$v2486\); 
          default_zero(\$v2379\); default_zero(\$v2139\); default_zero(cond); 
          default_zero(\$v177\); default_zero(\$v2037\); 
          default_zero(\$v251\); default_zero(\$v2381\); 
          default_zero(\$v2516\); default_zero(\$v2501\); 
          rdy <= "1";
          rdy1874 := "0";
          \state\ <= compute1875;
          state_var2552 <= compute2415;
          state_var2551 <= compute2412;
          state_var2550 <= compute2407;
          state_var2549 <= compute1922;
          
        else if run = '1' then
          case \state\ is
          when \$127_copy_args_to_heap544\ =>
            \$v1884\ := eclat_eq(\$127_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1884\(0) = '1' then
              \state\ <= \$127_copy_args_to_heap544\;
            else
              \$v1883\ := \$arr1869_ptr_take\;
              if \$v1883\(0) = '1' then
                \state\ <= q_wait1882;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$127_copy_args_to_heap544_arg\(32 to 63) & \$127_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                \state\ <= pause_getI1880;
              end if;
            end if;
          when \$128_pow568\ =>
            \$v1885\ := eclat_eq(\$128_pow568_arg\(32 to 63) & "00000000000000000000000000000000");
            if \$v1885\(0) = '1' then
              \state\ <= \$128_pow568\;
            else
              \$128_pow568_arg\ := \$128_pow568_arg\(0 to 31) & eclat_sub(\$128_pow568_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$128_pow568_arg\(64 to 95) & \$128_pow568_arg\(0 to 31));
              \state\ <= \$128_pow568\;
            end if;
          when \$129_div569\ =>
            \$v1894\ := eclat_eq(\$129_div569_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1894\(0) = '1' then
              \state\ <= \$129_div569\;
            else
              \$v1893\ := \$arr1869_ptr_take\;
              if \$v1893\(0) = '1' then
                \state\ <= q_wait1892;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$129_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$129_div569_arg\(0 to 31))));
                \state\ <= pause_getI1890;
              end if;
            end if;
          when \$130_mul570\ =>
            \$v1902\ := eclat_eq(\$130_mul570_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1902\(0) = '1' then
              \state\ <= \$130_mul570\;
            else
              \$v1901\ := \$arr1869_ptr_take\;
              if \$v1901\(0) = '1' then
                \state\ <= q_wait1900;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_mul570_arg\(0 to 31))));
                \state\ <= pause_getI1898;
              end if;
            end if;
          when \$131_sub571\ =>
            \$v1910\ := eclat_eq(\$131_sub571_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1910\(0) = '1' then
              \state\ <= \$131_sub571\;
            else
              \$v1909\ := \$arr1869_ptr_take\;
              if \$v1909\(0) = '1' then
                \state\ <= q_wait1908;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_sub571_arg\(0 to 31))));
                \state\ <= pause_getI1906;
              end if;
            end if;
          when \$132_add572\ =>
            \$v1918\ := eclat_eq(\$132_add572_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1918\(0) = '1' then
              \state\ <= \$132_add572\;
            else
              \$v1917\ := \$arr1869_ptr_take\;
              if \$v1917\(0) = '1' then
                \state\ <= q_wait1916;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_add572_arg\(0 to 31))));
                \state\ <= pause_getI1914;
              end if;
            end if;
          when \$615_forever5741837\ =>
            \state\ <= \$615_forever5741837\;
          when \$640_forever5741836\ =>
            \state\ <= \$640_forever5741836\;
          when \$665_forever5741835\ =>
            \state\ <= \$665_forever5741835\;
          when \$689_forever5741833\ =>
            \state\ <= \$689_forever5741833\;
          when \$698_forever5741834\ =>
            \state\ <= \$698_forever5741834\;
          when pause_getI1880 =>
            \state\ <= pause_getII1881;
          when pause_getI1890 =>
            \state\ <= pause_getII1891;
          when pause_getI1898 =>
            \state\ <= pause_getII1899;
          when pause_getI1906 =>
            \state\ <= pause_getII1907;
          when pause_getI1914 =>
            \state\ <= pause_getII1915;
          when pause_getII1881 =>
            \$arr1869_ptr_take\(0) := '0';
            \$726\ := \$arr1869_value\;
            \$v1879\ := \$arr1868_ptr_take\;
            if \$v1879\(0) = '1' then
              \state\ <= q_wait1878;
            else
              \$arr1868_ptr_take\(0) := '1';
              \$arr1868_ptr_write\ <= to_integer(unsigned(\$127_copy_args_to_heap544_arg\(64 to 95)));
              \$arr1868_write_request\ <= '1';
              \$arr1868_write\ <= \$726\;
              \state\ <= pause_setI1876;
            end if;
          when pause_getII1891 =>
            \$arr1869_ptr_take\(0) := '0';
            \$693\ := \$arr1869_value\;
            \$v1888\ := \$693\;
            \$v1889\ := \$v1888\(0 to 3);
            \$v1887\ := \$v1888\(4 to 67);
            case \$v1889\ is
            when "0001" =>
              \$694_a\ := \$v1887\(0 to 31);
              \$680_divisor\ := \$694_a\;
              \$v1886\ := eclat_eq(\$680_divisor\ & "00000000000000000000000000000000");
              if \$v1886\(0) = '1' then
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("Division par zero"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$689_forever5741833\;
              else
                \$129_div569_arg\ := eclat_sub(\$129_div569_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$129_div569_arg\(32 to 63) & \$680_divisor\) & \$129_div569_arg\(64 to 95);
                \state\ <= \$129_div569\;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$698_forever5741834\;
            end case;
          when pause_getII1899 =>
            \$arr1869_ptr_take\(0) := '0';
            \$655_v\ := \$arr1869_value\;
            \$v1896\ := \$655_v\;
            \$v1897\ := \$v1896\(0 to 3);
            \$v1895\ := \$v1896\(4 to 67);
            case \$v1897\ is
            when "0001" =>
              \$661_a\ := \$v1895\(0 to 31);
              \$656_int_value\ := \$661_a\;
              \$130_mul570_arg\ := eclat_sub(\$130_mul570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$130_mul570_arg\(32 to 63) & \$656_int_value\) & \$130_mul570_arg\(64 to 95);
              \state\ <= \$130_mul570\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$665_forever5741835\;
            end case;
          when pause_getII1907 =>
            \$arr1869_ptr_take\(0) := '0';
            \$630_v\ := \$arr1869_value\;
            \$v1904\ := \$630_v\;
            \$v1905\ := \$v1904\(0 to 3);
            \$v1903\ := \$v1904\(4 to 67);
            case \$v1905\ is
            when "0001" =>
              \$636_a\ := \$v1903\(0 to 31);
              \$631_int_value\ := \$636_a\;
              \$131_sub571_arg\ := eclat_sub(\$131_sub571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$131_sub571_arg\(32 to 63) & \$631_int_value\) & \$131_sub571_arg\(64 to 95);
              \state\ <= \$131_sub571\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$640_forever5741836\;
            end case;
          when pause_getII1915 =>
            \$arr1869_ptr_take\(0) := '0';
            \$605_v\ := \$arr1869_value\;
            \$v1912\ := \$605_v\;
            \$v1913\ := \$v1912\(0 to 3);
            \$v1911\ := \$v1912\(4 to 67);
            case \$v1913\ is
            when "0001" =>
              \$611_a\ := \$v1911\(0 to 31);
              \$606_int_value\ := \$611_a\;
              \$132_add572_arg\ := eclat_sub(\$132_add572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$132_add572_arg\(32 to 63) & \$606_int_value\) & \$132_add572_arg\(64 to 95);
              \state\ <= \$132_add572\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$615_forever5741837\;
            end case;
          when pause_setI1876 =>
            \$arr1868_write_request\ <= '0';
            \state\ <= pause_setII1877;
          when pause_setII1877 =>
            \$arr1868_ptr_take\(0) := '0';
            \$127_copy_args_to_heap544_arg\ := eclat_sub(\$127_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$127_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$127_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
            \state\ <= \$127_copy_args_to_heap544\;
          when q_wait1878 =>
            \$v1879\ := \$arr1868_ptr_take\;
            if \$v1879\(0) = '1' then
              \state\ <= q_wait1878;
            else
              \$arr1868_ptr_take\(0) := '1';
              \$arr1868_ptr_write\ <= to_integer(unsigned(\$127_copy_args_to_heap544_arg\(64 to 95)));
              \$arr1868_write_request\ <= '1';
              \$arr1868_write\ <= \$726\;
              \state\ <= pause_setI1876;
            end if;
          when q_wait1882 =>
            \$v1883\ := \$arr1869_ptr_take\;
            if \$v1883\(0) = '1' then
              \state\ <= q_wait1882;
            else
              \$arr1869_ptr_take\(0) := '1';
              \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$127_copy_args_to_heap544_arg\(32 to 63) & \$127_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI1880;
            end if;
          when q_wait1892 =>
            \$v1893\ := \$arr1869_ptr_take\;
            if \$v1893\(0) = '1' then
              \state\ <= q_wait1892;
            else
              \$arr1869_ptr_take\(0) := '1';
              \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$129_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$129_div569_arg\(0 to 31))));
              \state\ <= pause_getI1890;
            end if;
          when q_wait1900 =>
            \$v1901\ := \$arr1869_ptr_take\;
            if \$v1901\(0) = '1' then
              \state\ <= q_wait1900;
            else
              \$arr1869_ptr_take\(0) := '1';
              \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_mul570_arg\(0 to 31))));
              \state\ <= pause_getI1898;
            end if;
          when q_wait1908 =>
            \$v1909\ := \$arr1869_ptr_take\;
            if \$v1909\(0) = '1' then
              \state\ <= q_wait1908;
            else
              \$arr1869_ptr_take\(0) := '1';
              \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_sub571_arg\(0 to 31))));
              \state\ <= pause_getI1906;
            end if;
          when q_wait1916 =>
            \$v1917\ := \$arr1869_ptr_take\;
            if \$v1917\(0) = '1' then
              \state\ <= q_wait1916;
            else
              \$arr1869_ptr_take\(0) := '1';
              \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_add572_arg\(0 to 31))));
              \state\ <= pause_getI1914;
            end if;
          when compute1875 =>
            rdy1874 := eclat_false;
            case state_var2551 is
            when compute2412 =>
              rdy2411 := eclat_false;
              \$v2546\ := \$395\;
              if \$v2546\(0) = '1' then
                result2410 := eclat_true;
                rdy2411 := eclat_true;
                state_var2551 <= compute2412;
              else
                case state_var2552 is
                when \$400_copy_args_to_heap544\ =>
                  \$v2424\ := eclat_eq(\$400_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2424\(0) = '1' then
                    state_var2552 <= \$400_copy_args_to_heap544\;
                  else
                    \$v2423\ := \$arr1869_ptr_take\;
                    if \$v2423\(0) = '1' then
                      state_var2552 <= q_wait2422;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$400_copy_args_to_heap544_arg\(32 to 63) & \$400_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                      state_var2552 <= pause_getI2420;
                    end if;
                  end if;
                when \$401_pow568\ =>
                  \$v2425\ := eclat_eq(\$401_pow568_arg\(32 to 63) & "00000000000000000000000000000000");
                  if \$v2425\(0) = '1' then
                    state_var2552 <= \$401_pow568\;
                  else
                    \$401_pow568_arg\ := \$401_pow568_arg\(0 to 31) & eclat_sub(\$401_pow568_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$401_pow568_arg\(64 to 95) & \$401_pow568_arg\(0 to 31));
                    state_var2552 <= \$401_pow568\;
                  end if;
                when \$402_div569\ =>
                  \$v2434\ := eclat_eq(\$402_div569_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2434\(0) = '1' then
                    state_var2552 <= \$402_div569\;
                  else
                    \$v2433\ := \$arr1869_ptr_take\;
                    if \$v2433\(0) = '1' then
                      state_var2552 <= q_wait2432;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$402_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$402_div569_arg\(0 to 31))));
                      state_var2552 <= pause_getI2430;
                    end if;
                  end if;
                when \$403_mul570\ =>
                  \$v2442\ := eclat_eq(\$403_mul570_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2442\(0) = '1' then
                    state_var2552 <= \$403_mul570\;
                  else
                    \$v2441\ := \$arr1869_ptr_take\;
                    if \$v2441\(0) = '1' then
                      state_var2552 <= q_wait2440;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$403_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$403_mul570_arg\(0 to 31))));
                      state_var2552 <= pause_getI2438;
                    end if;
                  end if;
                when \$404_sub571\ =>
                  \$v2450\ := eclat_eq(\$404_sub571_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2450\(0) = '1' then
                    state_var2552 <= \$404_sub571\;
                  else
                    \$v2449\ := \$arr1869_ptr_take\;
                    if \$v2449\(0) = '1' then
                      state_var2552 <= q_wait2448;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$404_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$404_sub571_arg\(0 to 31))));
                      state_var2552 <= pause_getI2446;
                    end if;
                  end if;
                when \$405_add572\ =>
                  \$v2458\ := eclat_eq(\$405_add572_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2458\(0) = '1' then
                    state_var2552 <= \$405_add572\;
                  else
                    \$v2457\ := \$arr1869_ptr_take\;
                    if \$v2457\(0) = '1' then
                      state_var2552 <= q_wait2456;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$405_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$405_add572_arg\(0 to 31))));
                      state_var2552 <= pause_getI2454;
                    end if;
                  end if;
                when \$462_forever5741867\ =>
                  state_var2552 <= \$466_forever5741861\;
                when \$466_forever5741861\ =>
                  state_var2552 <= \$466_forever5741861\;
                when \$491_forever5741866\ =>
                  state_var2552 <= \$495_forever5741861\;
                when \$495_forever5741861\ =>
                  state_var2552 <= \$495_forever5741861\;
                when \$520_forever5741865\ =>
                  state_var2552 <= \$524_forever5741861\;
                when \$524_forever5741861\ =>
                  state_var2552 <= \$524_forever5741861\;
                when \$548_forever5741863\ =>
                  state_var2552 <= \$552_forever5741861\;
                when \$552_forever5741861\ =>
                  state_var2552 <= \$552_forever5741861\;
                when \$561_forever5741864\ =>
                  state_var2552 <= \$565_forever5741861\;
                when \$565_forever5741861\ =>
                  state_var2552 <= \$565_forever5741861\;
                when pause_getI2420 =>
                  state_var2552 <= pause_getII2421;
                when pause_getI2430 =>
                  state_var2552 <= pause_getII2431;
                when pause_getI2438 =>
                  state_var2552 <= pause_getII2439;
                when pause_getI2446 =>
                  state_var2552 <= pause_getII2447;
                when pause_getI2454 =>
                  state_var2552 <= pause_getII2455;
                when pause_getII2421 =>
                  \$arr1869_ptr_take\(0) := '0';
                  \$593\ := \$arr1869_value\;
                  \$v2419\ := \$arr1868_ptr_take\;
                  if \$v2419\(0) = '1' then
                    state_var2552 <= q_wait2418;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr_write\ <= to_integer(unsigned(\$400_copy_args_to_heap544_arg\(64 to 95)));
                    \$arr1868_write_request\ <= '1';
                    \$arr1868_write\ <= \$593\;
                    state_var2552 <= pause_setI2416;
                  end if;
                when pause_getII2431 =>
                  \$arr1869_ptr_take\(0) := '0';
                  \$556\ := \$arr1869_value\;
                  \$v2428\ := \$556\;
                  \$v2429\ := \$v2428\(0 to 3);
                  \$v2427\ := \$v2428\(4 to 67);
                  case \$v2429\ is
                  when "0001" =>
                    \$557_a\ := \$v2427\(0 to 31);
                    \$539_divisor\ := \$557_a\;
                    \$v2426\ := eclat_eq(\$539_divisor\ & "00000000000000000000000000000000");
                    if \$v2426\(0) = '1' then
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("Division par zero"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var2552 <= \$548_forever5741863\;
                    else
                      \$402_div569_arg\ := eclat_sub(\$402_div569_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$402_div569_arg\(32 to 63) & \$539_divisor\) & \$402_div569_arg\(64 to 95);
                      state_var2552 <= \$402_div569\;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2552 <= \$561_forever5741864\;
                  end case;
                when pause_getII2439 =>
                  \$arr1869_ptr_take\(0) := '0';
                  \$510_v\ := \$arr1869_value\;
                  \$v2436\ := \$510_v\;
                  \$v2437\ := \$v2436\(0 to 3);
                  \$v2435\ := \$v2436\(4 to 67);
                  case \$v2437\ is
                  when "0001" =>
                    \$516_a\ := \$v2435\(0 to 31);
                    \$511_int_value\ := \$516_a\;
                    \$403_mul570_arg\ := eclat_sub(\$403_mul570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$403_mul570_arg\(32 to 63) & \$511_int_value\) & \$403_mul570_arg\(64 to 95);
                    state_var2552 <= \$403_mul570\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2552 <= \$520_forever5741865\;
                  end case;
                when pause_getII2447 =>
                  \$arr1869_ptr_take\(0) := '0';
                  \$481_v\ := \$arr1869_value\;
                  \$v2444\ := \$481_v\;
                  \$v2445\ := \$v2444\(0 to 3);
                  \$v2443\ := \$v2444\(4 to 67);
                  case \$v2445\ is
                  when "0001" =>
                    \$487_a\ := \$v2443\(0 to 31);
                    \$482_int_value\ := \$487_a\;
                    \$404_sub571_arg\ := eclat_sub(\$404_sub571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$404_sub571_arg\(32 to 63) & \$482_int_value\) & \$404_sub571_arg\(64 to 95);
                    state_var2552 <= \$404_sub571\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2552 <= \$491_forever5741866\;
                  end case;
                when pause_getII2455 =>
                  \$arr1869_ptr_take\(0) := '0';
                  \$452_v\ := \$arr1869_value\;
                  \$v2452\ := \$452_v\;
                  \$v2453\ := \$v2452\(0 to 3);
                  \$v2451\ := \$v2452\(4 to 67);
                  case \$v2453\ is
                  when "0001" =>
                    \$458_a\ := \$v2451\(0 to 31);
                    \$453_int_value\ := \$458_a\;
                    \$405_add572_arg\ := eclat_sub(\$405_add572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$405_add572_arg\(32 to 63) & \$453_int_value\) & \$405_add572_arg\(64 to 95);
                    state_var2552 <= \$405_add572\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2552 <= \$462_forever5741867\;
                  end case;
                when pause_setI2416 =>
                  \$arr1868_write_request\ <= '0';
                  state_var2552 <= pause_setII2417;
                when pause_setI2460 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2461;
                when pause_setI2465 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2466;
                when pause_setI2470 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2471;
                when pause_setI2476 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2477;
                when pause_setI2482 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2483;
                when pause_setI2487 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2488;
                when pause_setI2492 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2493;
                when pause_setI2497 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2498;
                when pause_setI2503 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2504;
                when pause_setI2508 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2509;
                when pause_setI2513 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2514;
                when pause_setI2520 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2521;
                when pause_setI2525 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2526;
                when pause_setI2530 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2531;
                when pause_setI2535 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2536;
                when pause_setI2540 =>
                  \$arr1871_write_request\ <= '0';
                  state_var2552 <= pause_setII2541;
                when pause_setII2417 =>
                  \$arr1868_ptr_take\(0) := '0';
                  \$400_copy_args_to_heap544_arg\ := eclat_sub(\$400_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$400_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$400_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2552 <= \$400_copy_args_to_heap544\;
                when pause_setII2461 =>
                  \$arr1871_ptr_take\(0) := '0';
                  result2413 := eclat_unit;
                  rdy2414 := eclat_true;
                  state_var2552 <= compute2415;
                when pause_setII2466 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2463\ := \$arr1871_ptr_take\;
                  if \$v2463\(0) = '1' then
                    state_var2552 <= q_wait2462;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2459\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 15;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0111" & \$v2459\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2460;
                  end if;
                when pause_setII2471 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2468\ := \$arr1871_ptr_take\;
                  if \$v2468\(0) = '1' then
                    state_var2552 <= q_wait2467;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2464\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 14;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1000" & \$v2464\&X"000000000";
                    state_var2552 <= pause_setI2465;
                  end if;
                when pause_setII2477 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2473\ := \$arr1871_ptr_take\;
                  if \$v2473\(0) = '1' then
                    state_var2552 <= q_wait2472;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2469\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 13;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0010" & \$v2469\&X"000000000";
                    state_var2552 <= pause_setI2470;
                  end if;
                when pause_setII2483 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2479\ := \$arr1871_ptr_take\;
                  if \$v2479\(0) = '1' then
                    state_var2552 <= q_wait2478;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2474\ := "00000000000000000000000000000001";
                    \$v2475\ := "0001" & \$v2474\&X"00000000";
                    \$arr1871_ptr_write\ <= 12;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2475\;
                    state_var2552 <= pause_setI2476;
                  end if;
                when pause_setII2488 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2485\ := \$arr1871_ptr_take\;
                  if \$v2485\(0) = '1' then
                    state_var2552 <= q_wait2484;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2480\ := "00000000000000000000000000000010";
                    \$v2481\ := "0001" & \$v2480\&X"00000000";
                    \$arr1871_ptr_write\ <= 11;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2481\;
                    state_var2552 <= pause_setI2482;
                  end if;
                when pause_setII2493 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2490\ := \$arr1871_ptr_take\;
                  if \$v2490\(0) = '1' then
                    state_var2552 <= q_wait2489;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2486\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 10;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0001" & \$v2486\&X"000000000";
                    state_var2552 <= pause_setI2487;
                  end if;
                when pause_setII2498 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2495\ := \$arr1871_ptr_take\;
                  if \$v2495\(0) = '1' then
                    state_var2552 <= q_wait2494;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2491\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 9;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0110" & \$v2491\&X"000000000";
                    state_var2552 <= pause_setI2492;
                  end if;
                when pause_setII2504 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2500\ := \$arr1871_ptr_take\;
                  if \$v2500\(0) = '1' then
                    state_var2552 <= q_wait2499;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2496\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 8;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1001" & \$v2496\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2497;
                  end if;
                when pause_setII2509 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2506\ := \$arr1871_ptr_take\;
                  if \$v2506\(0) = '1' then
                    state_var2552 <= q_wait2505;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2501\ := eclat_unit;
                    \$v2502\ := "0010" & \$v2501\&"000"& X"000000000000000";
                    \$arr1871_ptr_write\ <= 7;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2502\;
                    state_var2552 <= pause_setI2503;
                  end if;
                when pause_setII2514 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2511\ := \$arr1871_ptr_take\;
                  if \$v2511\(0) = '1' then
                    state_var2552 <= q_wait2510;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2507\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 6;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1001" & \$v2507\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2508;
                  end if;
                when pause_setII2521 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2516\ := \$arr1871_ptr_take\;
                  if \$v2516\(0) = '1' then
                    state_var2552 <= q_wait2515;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2512\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 5;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1000" & \$v2512\&X"000000000";
                    state_var2552 <= pause_setI2513;
                  end if;
                when pause_setII2526 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2523\ := \$arr1871_ptr_take\;
                  if \$v2523\(0) = '1' then
                    state_var2552 <= q_wait2522;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2517\ := eclat_unit;
                    \$v2518\ := "0000" & \$v2517\;
                    \$v2519\ := "0011" & \$v2518\&"000"& X"00000000000000";
                    \$arr1871_ptr_write\ <= 4;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2519\;
                    state_var2552 <= pause_setI2520;
                  end if;
                when pause_setII2531 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2528\ := \$arr1871_ptr_take\;
                  if \$v2528\(0) = '1' then
                    state_var2552 <= q_wait2527;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2524\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 3;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0100" & \$v2524\&X"000000000";
                    state_var2552 <= pause_setI2525;
                  end if;
                when pause_setII2536 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2533\ := \$arr1871_ptr_take\;
                  if \$v2533\(0) = '1' then
                    state_var2552 <= q_wait2532;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2529\ := "00000000000000000000000000000001";
                    \$arr1871_ptr_write\ <= 2;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0100" & \$v2529\&X"000000000";
                    state_var2552 <= pause_setI2530;
                  end if;
                when pause_setII2541 =>
                  \$arr1871_ptr_take\(0) := '0';
                  \$v2538\ := \$arr1871_ptr_take\;
                  if \$v2538\(0) = '1' then
                    state_var2552 <= q_wait2537;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2534\ := "00000000000000000000000000001001";
                    \$arr1871_ptr_write\ <= 1;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1010" & \$v2534\&X"000000000";
                    state_var2552 <= pause_setI2535;
                  end if;
                when q_wait2418 =>
                  \$v2419\ := \$arr1868_ptr_take\;
                  if \$v2419\(0) = '1' then
                    state_var2552 <= q_wait2418;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr_write\ <= to_integer(unsigned(\$400_copy_args_to_heap544_arg\(64 to 95)));
                    \$arr1868_write_request\ <= '1';
                    \$arr1868_write\ <= \$593\;
                    state_var2552 <= pause_setI2416;
                  end if;
                when q_wait2422 =>
                  \$v2423\ := \$arr1869_ptr_take\;
                  if \$v2423\(0) = '1' then
                    state_var2552 <= q_wait2422;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$400_copy_args_to_heap544_arg\(32 to 63) & \$400_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var2552 <= pause_getI2420;
                  end if;
                when q_wait2432 =>
                  \$v2433\ := \$arr1869_ptr_take\;
                  if \$v2433\(0) = '1' then
                    state_var2552 <= q_wait2432;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$402_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$402_div569_arg\(0 to 31))));
                    state_var2552 <= pause_getI2430;
                  end if;
                when q_wait2440 =>
                  \$v2441\ := \$arr1869_ptr_take\;
                  if \$v2441\(0) = '1' then
                    state_var2552 <= q_wait2440;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$403_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$403_mul570_arg\(0 to 31))));
                    state_var2552 <= pause_getI2438;
                  end if;
                when q_wait2448 =>
                  \$v2449\ := \$arr1869_ptr_take\;
                  if \$v2449\(0) = '1' then
                    state_var2552 <= q_wait2448;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$404_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$404_sub571_arg\(0 to 31))));
                    state_var2552 <= pause_getI2446;
                  end if;
                when q_wait2456 =>
                  \$v2457\ := \$arr1869_ptr_take\;
                  if \$v2457\(0) = '1' then
                    state_var2552 <= q_wait2456;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$405_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$405_add572_arg\(0 to 31))));
                    state_var2552 <= pause_getI2454;
                  end if;
                when q_wait2462 =>
                  \$v2463\ := \$arr1871_ptr_take\;
                  if \$v2463\(0) = '1' then
                    state_var2552 <= q_wait2462;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2459\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 15;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0111" & \$v2459\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2460;
                  end if;
                when q_wait2467 =>
                  \$v2468\ := \$arr1871_ptr_take\;
                  if \$v2468\(0) = '1' then
                    state_var2552 <= q_wait2467;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2464\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 14;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1000" & \$v2464\&X"000000000";
                    state_var2552 <= pause_setI2465;
                  end if;
                when q_wait2472 =>
                  \$v2473\ := \$arr1871_ptr_take\;
                  if \$v2473\(0) = '1' then
                    state_var2552 <= q_wait2472;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2469\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 13;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0010" & \$v2469\&X"000000000";
                    state_var2552 <= pause_setI2470;
                  end if;
                when q_wait2478 =>
                  \$v2479\ := \$arr1871_ptr_take\;
                  if \$v2479\(0) = '1' then
                    state_var2552 <= q_wait2478;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2474\ := "00000000000000000000000000000001";
                    \$v2475\ := "0001" & \$v2474\&X"00000000";
                    \$arr1871_ptr_write\ <= 12;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2475\;
                    state_var2552 <= pause_setI2476;
                  end if;
                when q_wait2484 =>
                  \$v2485\ := \$arr1871_ptr_take\;
                  if \$v2485\(0) = '1' then
                    state_var2552 <= q_wait2484;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2480\ := "00000000000000000000000000000010";
                    \$v2481\ := "0001" & \$v2480\&X"00000000";
                    \$arr1871_ptr_write\ <= 11;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2481\;
                    state_var2552 <= pause_setI2482;
                  end if;
                when q_wait2489 =>
                  \$v2490\ := \$arr1871_ptr_take\;
                  if \$v2490\(0) = '1' then
                    state_var2552 <= q_wait2489;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2486\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 10;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0001" & \$v2486\&X"000000000";
                    state_var2552 <= pause_setI2487;
                  end if;
                when q_wait2494 =>
                  \$v2495\ := \$arr1871_ptr_take\;
                  if \$v2495\(0) = '1' then
                    state_var2552 <= q_wait2494;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2491\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 9;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0110" & \$v2491\&X"000000000";
                    state_var2552 <= pause_setI2492;
                  end if;
                when q_wait2499 =>
                  \$v2500\ := \$arr1871_ptr_take\;
                  if \$v2500\(0) = '1' then
                    state_var2552 <= q_wait2499;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2496\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 8;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1001" & \$v2496\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2497;
                  end if;
                when q_wait2505 =>
                  \$v2506\ := \$arr1871_ptr_take\;
                  if \$v2506\(0) = '1' then
                    state_var2552 <= q_wait2505;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2501\ := eclat_unit;
                    \$v2502\ := "0010" & \$v2501\&"000"& X"000000000000000";
                    \$arr1871_ptr_write\ <= 7;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2502\;
                    state_var2552 <= pause_setI2503;
                  end if;
                when q_wait2510 =>
                  \$v2511\ := \$arr1871_ptr_take\;
                  if \$v2511\(0) = '1' then
                    state_var2552 <= q_wait2510;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2507\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 6;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1001" & \$v2507\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2508;
                  end if;
                when q_wait2515 =>
                  \$v2516\ := \$arr1871_ptr_take\;
                  if \$v2516\(0) = '1' then
                    state_var2552 <= q_wait2515;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2512\ := "00000000000000000000000000000010";
                    \$arr1871_ptr_write\ <= 5;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1000" & \$v2512\&X"000000000";
                    state_var2552 <= pause_setI2513;
                  end if;
                when q_wait2522 =>
                  \$v2523\ := \$arr1871_ptr_take\;
                  if \$v2523\(0) = '1' then
                    state_var2552 <= q_wait2522;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2517\ := eclat_unit;
                    \$v2518\ := "0000" & \$v2517\;
                    \$v2519\ := "0011" & \$v2518\&"000"& X"00000000000000";
                    \$arr1871_ptr_write\ <= 4;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0101" & \$v2519\;
                    state_var2552 <= pause_setI2520;
                  end if;
                when q_wait2527 =>
                  \$v2528\ := \$arr1871_ptr_take\;
                  if \$v2528\(0) = '1' then
                    state_var2552 <= q_wait2527;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2524\ := "00000000000000000000000000000000";
                    \$arr1871_ptr_write\ <= 3;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0100" & \$v2524\&X"000000000";
                    state_var2552 <= pause_setI2525;
                  end if;
                when q_wait2532 =>
                  \$v2533\ := \$arr1871_ptr_take\;
                  if \$v2533\(0) = '1' then
                    state_var2552 <= q_wait2532;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2529\ := "00000000000000000000000000000001";
                    \$arr1871_ptr_write\ <= 2;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0100" & \$v2529\&X"000000000";
                    state_var2552 <= pause_setI2530;
                  end if;
                when q_wait2537 =>
                  \$v2538\ := \$arr1871_ptr_take\;
                  if \$v2538\(0) = '1' then
                    state_var2552 <= q_wait2537;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2534\ := "00000000000000000000000000001001";
                    \$arr1871_ptr_write\ <= 1;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "1010" & \$v2534\&X"000000000";
                    state_var2552 <= pause_setI2535;
                  end if;
                when q_wait2542 =>
                  \$v2543\ := \$arr1871_ptr_take\;
                  if \$v2543\(0) = '1' then
                    state_var2552 <= q_wait2542;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2539\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 0;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0000" & \$v2539\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2540;
                  end if;
                when compute2415 =>
                  rdy2414 := eclat_false;
                  \$v2543\ := \$arr1871_ptr_take\;
                  if \$v2543\(0) = '1' then
                    state_var2552 <= q_wait2542;
                  else
                    \$arr1871_ptr_take\(0) := '1';
                    \$v2539\ := eclat_unit;
                    \$arr1871_ptr_write\ <= 0;
                    \$arr1871_write_request\ <= '1';
                    \$arr1871_write\ <= "0000" & \$v2539\&"000"& X"0000000000000000";
                    state_var2552 <= pause_setI2540;
                  end if;
                end case;
                \$v2545\ := eclat_not(rdy2414);
                if \$v2545\(0) = '1' then
                  result2413 := eclat_unit;
                end if;
                \$397\ := result2413 & rdy2414;
                result2410 := ""&\$397\(1);
                rdy2411 := eclat_true;
                state_var2551 <= compute2412;
              end if;
            end case;
            \$v2548\ := eclat_not(rdy2411);
            if \$v2548\(0) = '1' then
              result2410 := eclat_false;
            end if;
            \$395\ := result2410;
            \$134_is_loaded\ := result2410;
            case state_var2550 is
            when compute2407 =>
              rdy2406 := eclat_false;
              result2405 := eclat_if(\$134_is_loaded\ & eclat_add(\$393\ & "00000000000000000000000000000001") & \$393\);
              rdy2406 := eclat_true;
              state_var2550 <= compute2407;
            end case;
            \$v2409\ := eclat_not(rdy2406);
            if \$v2409\(0) = '1' then
              result2405 := "00000000000000000000000000000000";
            end if;
            \$393\ := result2405;
            \$135_cy\ := result2405;
            case state_var2549 is
            when \$117_forever5731839\ =>
              state_var2549 <= \$117_forever5731839\;
            when \$117_forever5731846\ =>
              state_var2549 <= \$117_forever5731839\;
            when \$117_forever5731847\ =>
              state_var2549 <= \$117_forever5731839\;
            when \$117_forever5731848\ =>
              state_var2549 <= \$117_forever5731839\;
            when \$117_forever5731849\ =>
              state_var2549 <= \$117_forever5731839\;
            when \$120_forever5741838\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741850\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741851\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741852\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741853\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741854\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741855\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741856\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741857\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741858\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741859\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$120_forever5741860\ =>
              state_var2549 <= \$120_forever5741838\;
            when \$143_copy_args_to_heap544\ =>
              \$v1931\ := eclat_eq(\$143_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1931\(0) = '1' then
                \$143_copy_args_to_heap544_result\ := \$143_copy_args_to_heap544_arg\(32 to 63);
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(\$149_vm_run_code547_arg\(32 to 63));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2009\ := \$arr1868_ptr_take\;
                if \$v2009\(0) = '1' then
                  state_var2549 <= q_wait2008;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                  state_var2549 <= pause_getI2006;
                end if;
              else
                \$v1930\ := \$arr1869_ptr_take\;
                if \$v1930\(0) = '1' then
                  state_var2549 <= q_wait1929;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$143_copy_args_to_heap544_arg\(32 to 63) & \$143_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI1927;
                end if;
              end if;
            when \$144_pow568\ =>
              \$v1932\ := eclat_eq(\$144_pow568_arg\(32 to 63) & "00000000000000000000000000000000");
              if \$v1932\(0) = '1' then
                \$144_pow568_result\ := \$144_pow568_arg\(64 to 95);
                resultat := \$144_pow568_result\;
                \$v2138\ := \$arr1869_ptr_take\;
                if \$v2138\(0) = '1' then
                  state_var2549 <= q_wait2137;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2135;
                end if;
              else
                \$144_pow568_arg\ := \$144_pow568_arg\(0 to 31) & eclat_sub(\$144_pow568_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$144_pow568_arg\(64 to 95) & \$144_pow568_arg\(0 to 31));
                state_var2549 <= \$144_pow568\;
              end if;
            when \$145_div569\ =>
              \$v1941\ := eclat_eq(\$145_div569_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1941\(0) = '1' then
                \$145_div569_result\ := \$145_div569_arg\(32 to 63);
                resultat := \$145_div569_result\;
                \$v2157\ := \$arr1869_ptr_take\;
                if \$v2157\(0) = '1' then
                  state_var2549 <= q_wait2156;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2154;
                end if;
              else
                \$v1940\ := \$arr1869_ptr_take\;
                if \$v1940\(0) = '1' then
                  state_var2549 <= q_wait1939;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$145_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$145_div569_arg\(0 to 31))));
                  state_var2549 <= pause_getI1937;
                end if;
              end if;
            when \$146_mul570\ =>
              \$v1949\ := eclat_eq(\$146_mul570_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1949\(0) = '1' then
                \$146_mul570_result\ := \$146_mul570_arg\(32 to 63);
                resultat := \$146_mul570_result\;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2202\ := \$arr1869_ptr_take\;
                if \$v2202\(0) = '1' then
                  state_var2549 <= q_wait2201;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2199;
                end if;
              else
                \$v1948\ := \$arr1869_ptr_take\;
                if \$v1948\(0) = '1' then
                  state_var2549 <= q_wait1947;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_mul570_arg\(0 to 31))));
                  state_var2549 <= pause_getI1945;
                end if;
              end if;
            when \$147_sub571\ =>
              \$v1957\ := eclat_eq(\$147_sub571_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1957\(0) = '1' then
                \$147_sub571_result\ := \$147_sub571_arg\(32 to 63);
                resultat := \$147_sub571_result\;
                \$v2207\ := \$arr1869_ptr_take\;
                if \$v2207\(0) = '1' then
                  state_var2549 <= q_wait2206;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$v2203\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & \$v2203\&X"00000000";
                  state_var2549 <= pause_setI2204;
                end if;
              else
                \$v1956\ := \$arr1869_ptr_take\;
                if \$v1956\(0) = '1' then
                  state_var2549 <= q_wait1955;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_sub571_arg\(0 to 31))));
                  state_var2549 <= pause_getI1953;
                end if;
              end if;
            when \$148_add572\ =>
              \$v1965\ := eclat_eq(\$148_add572_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1965\(0) = '1' then
                \$148_add572_result\ := \$148_add572_arg\(32 to 63);
                resultat := \$148_add572_result\;
                \$v2252\ := \$arr1869_ptr_take\;
                if \$v2252\(0) = '1' then
                  state_var2549 <= q_wait2251;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2249;
                end if;
              else
                \$v1964\ := \$arr1869_ptr_take\;
                if \$v1964\(0) = '1' then
                  state_var2549 <= q_wait1963;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_add572_arg\(0 to 31))));
                  state_var2549 <= pause_getI1961;
                end if;
              end if;
            when \$149_vm_run_code547\ =>
              \$v2401\ := ""&\$149_vm_run_code547_arg\(294);
              if \$v2401\(0) = '1' then
                eclat_print_string(of_string("[sp:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(0 to 31));
                
                eclat_print_string(of_string("|env:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(32 to 63));
                
                eclat_print_string(of_string("|pc:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(64 to 95));
                
                eclat_print_string(of_string("|fp:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(96 to 127));
                
                eclat_print_string(of_string("]"));
                
                eclat_print_string(of_string("|gp:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(128 to 159));
                
                eclat_print_string(of_string("|hp:"));
                
                eclat_print_int(\$149_vm_run_code547_arg\(128 to 159));
                
                eclat_print_newline(eclat_unit);
                
                \$v2400\ := \$arr1871_ptr_take\;
                if \$v2400\(0) = '1' then
                  state_var2549 <= q_wait2399;
                else
                  \$arr1871_ptr_take\(0) := '1';
                  \$arr1871_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(64 to 95)));
                  state_var2549 <= pause_getI2397;
                end if;
              else
                \$v2400\ := \$arr1871_ptr_take\;
                if \$v2400\(0) = '1' then
                  state_var2549 <= q_wait2399;
                else
                  \$arr1871_ptr_take\(0) := '1';
                  \$arr1871_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(64 to 95)));
                  state_var2549 <= pause_getI2397;
                end if;
              end if;
            when \$208_forever5731845\ =>
              state_var2549 <= \$212_forever5731839\;
            when \$212_forever5731839\ =>
              state_var2549 <= \$212_forever5731839\;
            when \$258_forever5741844\ =>
              state_var2549 <= \$262_forever5741838\;
            when \$262_forever5741838\ =>
              state_var2549 <= \$262_forever5741838\;
            when \$287_forever5741843\ =>
              state_var2549 <= \$291_forever5741838\;
            when \$291_forever5741838\ =>
              state_var2549 <= \$291_forever5741838\;
            when \$316_forever5741842\ =>
              state_var2549 <= \$320_forever5741838\;
            when \$320_forever5741838\ =>
              state_var2549 <= \$320_forever5741838\;
            when \$344_forever5741840\ =>
              state_var2549 <= \$348_forever5741838\;
            when \$348_forever5741838\ =>
              state_var2549 <= \$348_forever5741838\;
            when \$357_forever5741841\ =>
              state_var2549 <= \$361_forever5741838\;
            when \$361_forever5741838\ =>
              state_var2549 <= \$361_forever5741838\;
            when pause_getI1927 =>
              state_var2549 <= pause_getII1928;
            when pause_getI1937 =>
              state_var2549 <= pause_getII1938;
            when pause_getI1945 =>
              state_var2549 <= pause_getII1946;
            when pause_getI1953 =>
              state_var2549 <= pause_getII1954;
            when pause_getI1961 =>
              state_var2549 <= pause_getII1962;
            when pause_getI1984 =>
              state_var2549 <= pause_getII1985;
            when pause_getI1995 =>
              state_var2549 <= pause_getII1996;
            when pause_getI2006 =>
              state_var2549 <= pause_getII2007;
            when pause_getI2017 =>
              state_var2549 <= pause_getII2018;
            when pause_getI2028 =>
              state_var2549 <= pause_getII2029;
            when pause_getI2039 =>
              state_var2549 <= pause_getII2040;
            when pause_getI2065 =>
              state_var2549 <= pause_getII2066;
            when pause_getI2069 =>
              state_var2549 <= pause_getII2070;
            when pause_getI2094 =>
              state_var2549 <= pause_getII2095;
            when pause_getI2105 =>
              state_var2549 <= pause_getII2106;
            when pause_getI2116 =>
              state_var2549 <= pause_getII2117;
            when pause_getI2123 =>
              state_var2549 <= pause_getII2124;
            when pause_getI2130 =>
              state_var2549 <= pause_getII2131;
            when pause_getI2142 =>
              state_var2549 <= pause_getII2143;
            when pause_getI2149 =>
              state_var2549 <= pause_getII2150;
            when pause_getI2161 =>
              state_var2549 <= pause_getII2162;
            when pause_getI2177 =>
              state_var2549 <= pause_getII2178;
            when pause_getI2188 =>
              state_var2549 <= pause_getII2189;
            when pause_getI2199 =>
              state_var2549 <= pause_getII2200;
            when pause_getI2215 =>
              state_var2549 <= pause_getII2216;
            when pause_getI2226 =>
              state_var2549 <= pause_getII2227;
            when pause_getI2237 =>
              state_var2549 <= pause_getII2238;
            when pause_getI2244 =>
              state_var2549 <= pause_getII2245;
            when pause_getI2260 =>
              state_var2549 <= pause_getII2261;
            when pause_getI2271 =>
              state_var2549 <= pause_getII2272;
            when pause_getI2282 =>
              state_var2549 <= pause_getII2283;
            when pause_getI2290 =>
              state_var2549 <= pause_getII2291;
            when pause_getI2303 =>
              state_var2549 <= pause_getII2304;
            when pause_getI2307 =>
              state_var2549 <= pause_getII2308;
            when pause_getI2314 =>
              state_var2549 <= pause_getII2315;
            when pause_getI2321 =>
              state_var2549 <= pause_getII2322;
            when pause_getI2329 =>
              state_var2549 <= pause_getII2330;
            when pause_getI2337 =>
              state_var2549 <= pause_getII2338;
            when pause_getI2348 =>
              state_var2549 <= pause_getII2349;
            when pause_getI2359 =>
              state_var2549 <= pause_getII2360;
            when pause_getI2367 =>
              state_var2549 <= pause_getII2368;
            when pause_getI2375 =>
              state_var2549 <= pause_getII2376;
            when pause_getI2386 =>
              state_var2549 <= pause_getII2387;
            when pause_getI2397 =>
              state_var2549 <= pause_getII2398;
            when pause_getII1928 =>
              \$arr1869_ptr_take\(0) := '0';
              \$389\ := \$arr1869_value\;
              \$v1926\ := \$arr1868_ptr_take\;
              if \$v1926\(0) = '1' then
                state_var2549 <= q_wait1925;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr_write\ <= to_integer(unsigned(\$143_copy_args_to_heap544_arg\(64 to 95)));
                \$arr1868_write_request\ <= '1';
                \$arr1868_write\ <= \$389\;
                state_var2549 <= pause_setI1923;
              end if;
            when pause_getII1938 =>
              \$arr1869_ptr_take\(0) := '0';
              \$352\ := \$arr1869_value\;
              \$v1935\ := \$352\;
              \$v1936\ := \$v1935\(0 to 3);
              \$v1934\ := \$v1935\(4 to 67);
              case \$v1936\ is
              when "0001" =>
                \$353_a\ := \$v1934\(0 to 31);
                \$335_divisor\ := \$353_a\;
                \$v1933\ := eclat_eq(\$335_divisor\ & "00000000000000000000000000000000");
                if \$v1933\(0) = '1' then
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("Division par zero"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2549 <= \$344_forever5741840\;
                else
                  \$145_div569_arg\ := eclat_sub(\$145_div569_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$145_div569_arg\(32 to 63) & \$335_divisor\) & \$145_div569_arg\(64 to 95);
                  state_var2549 <= \$145_div569\;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$357_forever5741841\;
              end case;
            when pause_getII1946 =>
              \$arr1869_ptr_take\(0) := '0';
              \$306_v\ := \$arr1869_value\;
              \$v1943\ := \$306_v\;
              \$v1944\ := \$v1943\(0 to 3);
              \$v1942\ := \$v1943\(4 to 67);
              case \$v1944\ is
              when "0001" =>
                \$312_a\ := \$v1942\(0 to 31);
                \$307_int_value\ := \$312_a\;
                \$146_mul570_arg\ := eclat_sub(\$146_mul570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$146_mul570_arg\(32 to 63) & \$307_int_value\) & \$146_mul570_arg\(64 to 95);
                state_var2549 <= \$146_mul570\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$316_forever5741842\;
              end case;
            when pause_getII1954 =>
              \$arr1869_ptr_take\(0) := '0';
              \$277_v\ := \$arr1869_value\;
              \$v1951\ := \$277_v\;
              \$v1952\ := \$v1951\(0 to 3);
              \$v1950\ := \$v1951\(4 to 67);
              case \$v1952\ is
              when "0001" =>
                \$283_a\ := \$v1950\(0 to 31);
                \$278_int_value\ := \$283_a\;
                \$147_sub571_arg\ := eclat_sub(\$147_sub571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$147_sub571_arg\(32 to 63) & \$278_int_value\) & \$147_sub571_arg\(64 to 95);
                state_var2549 <= \$147_sub571\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$287_forever5741843\;
              end case;
            when pause_getII1962 =>
              \$arr1869_ptr_take\(0) := '0';
              \$248_v\ := \$arr1869_value\;
              \$v1959\ := \$248_v\;
              \$v1960\ := \$v1959\(0 to 3);
              \$v1958\ := \$v1959\(4 to 67);
              case \$v1960\ is
              when "0001" =>
                \$254_a\ := \$v1958\(0 to 31);
                \$249_int_value\ := \$254_a\;
                \$148_add572_arg\ := eclat_sub(\$148_add572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$148_add572_arg\(32 to 63) & \$249_int_value\) & \$148_add572_arg\(64 to 95);
                state_var2549 <= \$148_add572\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$258_forever5741844\;
              end case;
            when pause_getII1985 =>
              \$arr1868_ptr_take\(0) := '0';
              \$v42\ := \$arr1868_value\;
              \$v1982\ := \$v42\;
              \$v1983\ := \$v1982\(0 to 3);
              \$v1977\ := \$v1982\(4 to 67);
              case \$v1983\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1976\ := \$arr1872_ptr_take\;
                if \$v1976\(0) = '1' then
                  state_var2549 <= q_wait1975;
                else
                  \$arr1872_ptr_take\(0) := '1';
                  \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                  \$arr1872_write_request\ <= '1';
                  \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                  state_var2549 <= pause_setI1973;
                end if;
              when "0011" =>
                \$113_p\ := \$v1977\(0 to 4);
                \$v1979\ := \$113_p\;
                \$v1980\ := \$v1979\(0 to 3);
                \$v1978\ := ""&\$v1979\(4);
                case \$v1980\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1976\ := \$arr1872_ptr_take\;
                if \$v1976\(0) = '1' then
                  state_var2549 <= q_wait1975;
                else
                  \$arr1872_ptr_take\(0) := '1';
                  \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                  \$arr1872_write_request\ <= '1';
                  \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                  state_var2549 <= pause_setI1973;
                end if;
              when "0001" =>
                \$114_n\ := \$v1977\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v1976\ := \$arr1872_ptr_take\;
                if \$v1976\(0) = '1' then
                  state_var2549 <= q_wait1975;
                else
                  \$arr1872_ptr_take\(0) := '1';
                  \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                  \$arr1872_write_request\ <= '1';
                  \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                  state_var2549 <= pause_setI1973;
                end if;
              when "0000" =>
                \$115_b\ := \$v1977\(0 to 0);
                \$v1981\ := \$115_b\;
                if \$v1981\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1976\ := \$arr1872_ptr_take\;
                  if \$v1976\(0) = '1' then
                    state_var2549 <= q_wait1975;
                  else
                    \$arr1872_ptr_take\(0) := '1';
                    \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                    \$arr1872_write_request\ <= '1';
                    \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                    state_var2549 <= pause_setI1973;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1996 =>
              \$arr1868_ptr_take\(0) := '0';
              \$v39\ := \$arr1868_value\;
              \$v1993\ := \$v39\;
              \$v1994\ := \$v1993\(0 to 3);
              \$v1988\ := \$v1993\(4 to 67);
              case \$v1994\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1987\ := \$arr1868_ptr_take\;
                if \$v1987\(0) = '1' then
                  state_var2549 <= q_wait1986;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI1984;
                end if;
              when "0011" =>
                \$113_p\ := \$v1988\(0 to 4);
                \$v1990\ := \$113_p\;
                \$v1991\ := \$v1990\(0 to 3);
                \$v1989\ := ""&\$v1990\(4);
                case \$v1991\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1987\ := \$arr1868_ptr_take\;
                if \$v1987\(0) = '1' then
                  state_var2549 <= q_wait1986;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI1984;
                end if;
              when "0001" =>
                \$114_n\ := \$v1988\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1987\ := \$arr1868_ptr_take\;
                if \$v1987\(0) = '1' then
                  state_var2549 <= q_wait1986;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI1984;
                end if;
              when "0000" =>
                \$115_b\ := \$v1988\(0 to 0);
                \$v1992\ := \$115_b\;
                if \$v1992\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1987\ := \$arr1868_ptr_take\;
                  if \$v1987\(0) = '1' then
                    state_var2549 <= q_wait1986;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI1984;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2007 =>
              \$arr1868_ptr_take\(0) := '0';
              \$v36\ := \$arr1868_value\;
              \$v2004\ := \$v36\;
              \$v2005\ := \$v2004\(0 to 3);
              \$v1999\ := \$v2004\(4 to 67);
              case \$v2005\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1998\ := \$arr1868_ptr_take\;
                if \$v1998\(0) = '1' then
                  state_var2549 <= q_wait1997;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI1995;
                end if;
              when "0011" =>
                \$113_p\ := \$v1999\(0 to 4);
                \$v2001\ := \$113_p\;
                \$v2002\ := \$v2001\(0 to 3);
                \$v2000\ := ""&\$v2001\(4);
                case \$v2002\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1998\ := \$arr1868_ptr_take\;
                if \$v1998\(0) = '1' then
                  state_var2549 <= q_wait1997;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI1995;
                end if;
              when "0001" =>
                \$114_n\ := \$v1999\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("heap["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1998\ := \$arr1868_ptr_take\;
                if \$v1998\(0) = '1' then
                  state_var2549 <= q_wait1997;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI1995;
                end if;
              when "0000" =>
                \$115_b\ := \$v1999\(0 to 0);
                \$v2003\ := \$115_b\;
                if \$v2003\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("heap["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1998\ := \$arr1868_ptr_take\;
                  if \$v1998\(0) = '1' then
                    state_var2549 <= q_wait1997;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI1995;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2018 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v33\ := \$arr1869_value\;
              \$v2015\ := \$v33\;
              \$v2016\ := \$v2015\(0 to 3);
              \$v2010\ := \$v2015\(4 to 67);
              case \$v2016\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                state_var2549 <= \$143_copy_args_to_heap544\;
              when "0011" =>
                \$113_p\ := \$v2010\(0 to 4);
                \$v2012\ := \$113_p\;
                \$v2013\ := \$v2012\(0 to 3);
                \$v2011\ := ""&\$v2012\(4);
                case \$v2013\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                state_var2549 <= \$143_copy_args_to_heap544\;
              when "0001" =>
                \$114_n\ := \$v2010\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                state_var2549 <= \$143_copy_args_to_heap544\;
              when "0000" =>
                \$115_b\ := \$v2010\(0 to 0);
                \$v2014\ := \$115_b\;
                if \$v2014\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$143_copy_args_to_heap544_arg\ := \$192_n\ & \$149_vm_run_code547_arg\(0 to 31) & eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001");
                  state_var2549 <= \$143_copy_args_to_heap544\;
                end if;
              when others =>
                
              end case;
            when pause_getII2029 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v26\ := \$arr1869_value\;
              \$v2026\ := \$v26\;
              \$v2027\ := \$v2026\(0 to 3);
              \$v2021\ := \$v2026\(4 to 67);
              case \$v2027\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2020\ := \$arr1869_ptr_take\;
                if \$v2020\(0) = '1' then
                  state_var2549 <= q_wait2019;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2017;
                end if;
              when "0011" =>
                \$113_p\ := \$v2021\(0 to 4);
                \$v2023\ := \$113_p\;
                \$v2024\ := \$v2023\(0 to 3);
                \$v2022\ := ""&\$v2023\(4);
                case \$v2024\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2020\ := \$arr1869_ptr_take\;
                if \$v2020\(0) = '1' then
                  state_var2549 <= q_wait2019;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2017;
                end if;
              when "0001" =>
                \$114_n\ := \$v2021\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2020\ := \$arr1869_ptr_take\;
                if \$v2020\(0) = '1' then
                  state_var2549 <= q_wait2019;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2017;
                end if;
              when "0000" =>
                \$115_b\ := \$v2021\(0 to 0);
                \$v2025\ := \$115_b\;
                if \$v2025\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2020\ := \$arr1869_ptr_take\;
                  if \$v2020\(0) = '1' then
                    state_var2549 <= q_wait2019;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2017;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2040 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v23\ := \$arr1869_value\;
              \$v2037\ := \$v23\;
              \$v2038\ := \$v2037\(0 to 3);
              \$v2032\ := \$v2037\(4 to 67);
              case \$v2038\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2031\ := \$arr1869_ptr_take\;
                if \$v2031\(0) = '1' then
                  state_var2549 <= q_wait2030;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2028;
                end if;
              when "0011" =>
                \$113_p\ := \$v2032\(0 to 4);
                \$v2034\ := \$113_p\;
                \$v2035\ := \$v2034\(0 to 3);
                \$v2033\ := ""&\$v2034\(4);
                case \$v2035\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2031\ := \$arr1869_ptr_take\;
                if \$v2031\(0) = '1' then
                  state_var2549 <= q_wait2030;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2028;
                end if;
              when "0001" =>
                \$114_n\ := \$v2032\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2031\ := \$arr1869_ptr_take\;
                if \$v2031\(0) = '1' then
                  state_var2549 <= q_wait2030;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2028;
                end if;
              when "0000" =>
                \$115_b\ := \$v2032\(0 to 0);
                \$v2036\ := \$115_b\;
                if \$v2036\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2031\ := \$arr1869_ptr_take\;
                  if \$v2031\(0) = '1' then
                    state_var2549 <= q_wait2030;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2028;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2066 =>
              \$arr1869_ptr_take\(0) := '0';
              second_value := \$arr1869_value\;
              \$v2063\ := first_value;
              \$v2064\ := \$v2063\(0 to 3);
              \$v2053\ := \$v2063\(4 to 67);
              case \$v2064\ is
              when "0010" =>
                \$v2055\ := second_value;
                \$v2056\ := \$v2055\(0 to 3);
                \$v2054\ := \$v2055\(4 to 67);
                case \$v2056\ is
                when "0010" =>
                  res := eclat_true;
                  \$v2052\ := \$arr1869_ptr_take\;
                  if \$v2052\(0) = '1' then
                    state_var2549 <= q_wait2051;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2049;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2549 <= \$117_forever5731847\;
                end case;
              when "0000" =>
                \$98_a1\ := \$v2053\(0 to 0);
                \$v2058\ := second_value;
                \$v2059\ := \$v2058\(0 to 3);
                \$v2057\ := \$v2058\(4 to 67);
                case \$v2059\ is
                when "0000" =>
                  b2 := \$v2057\(0 to 0);
                  res := eclat_if(\$98_a1\ & eclat_if(b2 & eclat_true & eclat_false) & 
                         eclat_if(b2 & eclat_false & eclat_true));
                  \$v2052\ := \$arr1869_ptr_take\;
                  if \$v2052\(0) = '1' then
                    state_var2549 <= q_wait2051;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2049;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2549 <= \$117_forever5731848\;
                end case;
              when "0001" =>
                \$99_a\ := \$v2053\(0 to 31);
                \$v2061\ := second_value;
                \$v2062\ := \$v2061\(0 to 3);
                \$v2060\ := \$v2061\(4 to 67);
                case \$v2062\ is
                when "0001" =>
                  b := \$v2060\(0 to 31);
                  res := eclat_eq(\$99_a\ & b);
                  \$v2052\ := \$arr1869_ptr_take\;
                  if \$v2052\(0) = '1' then
                    state_var2549 <= q_wait2051;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2049;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2549 <= \$117_forever5731849\;
                end case;
              when others =>
                eclat_print_string(of_string("il n'y a pas d'égalité possible \n"));
                
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$117_forever5731846\;
              end case;
            when pause_getII2070 =>
              \$arr1869_ptr_take\(0) := '0';
              first_value := \$arr1869_value\;
              \$v2068\ := \$arr1869_ptr_take\;
              if \$v2068\(0) = '1' then
                state_var2549 <= q_wait2067;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2549 <= pause_getI2065;
              end if;
            when pause_getII2095 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v81\ := \$arr1869_value\;
              \$v2092\ := \$v81\;
              \$v2093\ := \$v2092\(0 to 3);
              \$v2087\ := \$v2092\(4 to 67);
              case \$v2093\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2086\ := \$arr1869_ptr_take\;
                if \$v2086\(0) = '1' then
                  state_var2549 <= q_wait2085;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$v2082\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                  state_var2549 <= pause_setI2083;
                end if;
              when "0011" =>
                \$113_p\ := \$v2087\(0 to 4);
                \$v2089\ := \$113_p\;
                \$v2090\ := \$v2089\(0 to 3);
                \$v2088\ := ""&\$v2089\(4);
                case \$v2090\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2086\ := \$arr1869_ptr_take\;
                if \$v2086\(0) = '1' then
                  state_var2549 <= q_wait2085;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$v2082\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                  state_var2549 <= pause_setI2083;
                end if;
              when "0001" =>
                \$114_n\ := \$v2087\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v2086\ := \$arr1869_ptr_take\;
                if \$v2086\(0) = '1' then
                  state_var2549 <= q_wait2085;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$v2082\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                  state_var2549 <= pause_setI2083;
                end if;
              when "0000" =>
                \$115_b\ := \$v2087\(0 to 0);
                \$v2091\ := \$115_b\;
                if \$v2091\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2086\ := \$arr1869_ptr_take\;
                  if \$v2086\(0) = '1' then
                    state_var2549 <= q_wait2085;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$v2082\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                    state_var2549 <= pause_setI2083;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2106 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v78\ := \$arr1869_value\;
              \$v2103\ := \$v78\;
              \$v2104\ := \$v2103\(0 to 3);
              \$v2098\ := \$v2103\(4 to 67);
              case \$v2104\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2097\ := \$arr1869_ptr_take\;
                if \$v2097\(0) = '1' then
                  state_var2549 <= q_wait2096;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2094;
                end if;
              when "0011" =>
                \$113_p\ := \$v2098\(0 to 4);
                \$v2100\ := \$113_p\;
                \$v2101\ := \$v2100\(0 to 3);
                \$v2099\ := ""&\$v2100\(4);
                case \$v2101\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2097\ := \$arr1869_ptr_take\;
                if \$v2097\(0) = '1' then
                  state_var2549 <= q_wait2096;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2094;
                end if;
              when "0001" =>
                \$114_n\ := \$v2098\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2097\ := \$arr1869_ptr_take\;
                if \$v2097\(0) = '1' then
                  state_var2549 <= q_wait2096;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2094;
                end if;
              when "0000" =>
                \$115_b\ := \$v2098\(0 to 0);
                \$v2102\ := \$115_b\;
                if \$v2102\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2097\ := \$arr1869_ptr_take\;
                  if \$v2097\(0) = '1' then
                    state_var2549 <= q_wait2096;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2094;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2117 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v75\ := \$arr1869_value\;
              \$v2114\ := \$v75\;
              \$v2115\ := \$v2114\(0 to 3);
              \$v2109\ := \$v2114\(4 to 67);
              case \$v2115\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2108\ := \$arr1869_ptr_take\;
                if \$v2108\(0) = '1' then
                  state_var2549 <= q_wait2107;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI2105;
                end if;
              when "0011" =>
                \$113_p\ := \$v2109\(0 to 4);
                \$v2111\ := \$113_p\;
                \$v2112\ := \$v2111\(0 to 3);
                \$v2110\ := ""&\$v2111\(4);
                case \$v2112\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2108\ := \$arr1869_ptr_take\;
                if \$v2108\(0) = '1' then
                  state_var2549 <= q_wait2107;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI2105;
                end if;
              when "0001" =>
                \$114_n\ := \$v2109\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2108\ := \$arr1869_ptr_take\;
                if \$v2108\(0) = '1' then
                  state_var2549 <= q_wait2107;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI2105;
                end if;
              when "0000" =>
                \$115_b\ := \$v2109\(0 to 0);
                \$v2113\ := \$115_b\;
                if \$v2113\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2108\ := \$arr1869_ptr_take\;
                  if \$v2108\(0) = '1' then
                    state_var2549 <= q_wait2107;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2549 <= pause_getI2105;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2124 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v72\ := \$arr1869_value\;
              \$v2121\ := \$v72\;
              \$v2122\ := \$v2121\(0 to 3);
              \$v2120\ := \$v2121\(4 to 67);
              case \$v2122\ is
              when "0001" =>
                a := \$v2120\(0 to 31);
                scd_operand := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2119\ := \$arr1869_ptr_take\;
                if \$v2119\(0) = '1' then
                  state_var2549 <= q_wait2118;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                  state_var2549 <= pause_getI2116;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741851\;
              end case;
            when pause_getII2131 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v70\ := \$arr1869_value\;
              \$v2128\ := \$v70\;
              \$v2129\ := \$v2128\(0 to 3);
              \$v2127\ := \$v2128\(4 to 67);
              case \$v2129\ is
              when "0001" =>
                a := \$v2127\(0 to 31);
                fst_operand := a;
                \$v2126\ := \$arr1869_ptr_take\;
                if \$v2126\(0) = '1' then
                  state_var2549 <= q_wait2125;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI2123;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741852\;
              end case;
            when pause_getII2143 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v93\ := \$arr1869_value\;
              \$v2140\ := \$v93\;
              \$v2141\ := \$v2140\(0 to 3);
              \$v2139\ := \$v2140\(4 to 67);
              case \$v2141\ is
              when "0001" =>
                a := \$v2139\(0 to 31);
                exponent := a;
                \$144_pow568_arg\ := base & exponent & "00000000000000000000000000000001";
                state_var2549 <= \$144_pow568\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741854\;
              end case;
            when pause_getII2150 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v91\ := \$arr1869_value\;
              \$v2147\ := \$v91\;
              \$v2148\ := \$v2147\(0 to 3);
              \$v2146\ := \$v2147\(4 to 67);
              case \$v2148\ is
              when "0001" =>
                a := \$v2146\(0 to 31);
                base := a;
                \$v2145\ := \$arr1869_ptr_take\;
                if \$v2145\(0) = '1' then
                  state_var2549 <= q_wait2144;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2549 <= pause_getI2142;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741855\;
              end case;
            when pause_getII2162 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v117\ := \$arr1869_value\;
              \$v2159\ := \$v117\;
              \$v2160\ := \$v2159\(0 to 3);
              \$v2158\ := \$v2159\(4 to 67);
              case \$v2160\ is
              when "0001" =>
                a := \$v2158\(0 to 31);
                debut := a;
                \$145_div569_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$145_div569\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741857\;
              end case;
            when pause_getII2178 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v149\ := \$arr1869_value\;
              \$v2175\ := \$v149\;
              \$v2176\ := \$v2175\(0 to 3);
              \$v2170\ := \$v2175\(4 to 67);
              case \$v2176\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2169\ := \$arr1869_ptr_take\;
                if \$v2169\(0) = '1' then
                  state_var2549 <= q_wait2168;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2166;
                end if;
              when "0011" =>
                \$113_p\ := \$v2170\(0 to 4);
                \$v2172\ := \$113_p\;
                \$v2173\ := \$v2172\(0 to 3);
                \$v2171\ := ""&\$v2172\(4);
                case \$v2173\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2169\ := \$arr1869_ptr_take\;
                if \$v2169\(0) = '1' then
                  state_var2549 <= q_wait2168;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2166;
                end if;
              when "0001" =>
                \$114_n\ := \$v2170\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v2169\ := \$arr1869_ptr_take\;
                if \$v2169\(0) = '1' then
                  state_var2549 <= q_wait2168;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0001" & resultat&X"00000000";
                  state_var2549 <= pause_setI2166;
                end if;
              when "0000" =>
                \$115_b\ := \$v2170\(0 to 0);
                \$v2174\ := \$115_b\;
                if \$v2174\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2169\ := \$arr1869_ptr_take\;
                  if \$v2169\(0) = '1' then
                    state_var2549 <= q_wait2168;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1869_write_request\ <= '1';
                    \$arr1869_write\ <= "0001" & resultat&X"00000000";
                    state_var2549 <= pause_setI2166;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2189 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v142\ := \$arr1869_value\;
              \$v2186\ := \$v142\;
              \$v2187\ := \$v2186\(0 to 3);
              \$v2181\ := \$v2186\(4 to 67);
              case \$v2187\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2180\ := \$arr1869_ptr_take\;
                if \$v2180\(0) = '1' then
                  state_var2549 <= q_wait2179;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2177;
                end if;
              when "0011" =>
                \$113_p\ := \$v2181\(0 to 4);
                \$v2183\ := \$113_p\;
                \$v2184\ := \$v2183\(0 to 3);
                \$v2182\ := ""&\$v2183\(4);
                case \$v2184\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2180\ := \$arr1869_ptr_take\;
                if \$v2180\(0) = '1' then
                  state_var2549 <= q_wait2179;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2177;
                end if;
              when "0001" =>
                \$114_n\ := \$v2181\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2180\ := \$arr1869_ptr_take\;
                if \$v2180\(0) = '1' then
                  state_var2549 <= q_wait2179;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2177;
                end if;
              when "0000" =>
                \$115_b\ := \$v2181\(0 to 0);
                \$v2185\ := \$115_b\;
                if \$v2185\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2180\ := \$arr1869_ptr_take\;
                  if \$v2180\(0) = '1' then
                    state_var2549 <= q_wait2179;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2177;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2200 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v139\ := \$arr1869_value\;
              \$v2197\ := \$v139\;
              \$v2198\ := \$v2197\(0 to 3);
              \$v2192\ := \$v2197\(4 to 67);
              case \$v2198\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2191\ := \$arr1869_ptr_take\;
                if \$v2191\(0) = '1' then
                  state_var2549 <= q_wait2190;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2188;
                end if;
              when "0011" =>
                \$113_p\ := \$v2192\(0 to 4);
                \$v2194\ := \$113_p\;
                \$v2195\ := \$v2194\(0 to 3);
                \$v2193\ := ""&\$v2194\(4);
                case \$v2195\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2191\ := \$arr1869_ptr_take\;
                if \$v2191\(0) = '1' then
                  state_var2549 <= q_wait2190;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2188;
                end if;
              when "0001" =>
                \$114_n\ := \$v2192\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2191\ := \$arr1869_ptr_take\;
                if \$v2191\(0) = '1' then
                  state_var2549 <= q_wait2190;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2188;
                end if;
              when "0000" =>
                \$115_b\ := \$v2192\(0 to 0);
                \$v2196\ := \$115_b\;
                if \$v2196\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2191\ := \$arr1869_ptr_take\;
                  if \$v2191\(0) = '1' then
                    state_var2549 <= q_wait2190;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2188;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2216 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v184\ := \$arr1869_value\;
              \$v2213\ := \$v184\;
              \$v2214\ := \$v2213\(0 to 3);
              \$v2208\ := \$v2213\(4 to 67);
              case \$v2214\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$147_sub571\;
              when "0011" =>
                \$113_p\ := \$v2208\(0 to 4);
                \$v2210\ := \$113_p\;
                \$v2211\ := \$v2210\(0 to 3);
                \$v2209\ := ""&\$v2210\(4);
                case \$v2211\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$147_sub571\;
              when "0001" =>
                \$114_n\ := \$v2208\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$147_sub571\;
              when "0000" =>
                \$115_b\ := \$v2208\(0 to 0);
                \$v2212\ := \$115_b\;
                if \$v2212\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub571_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$147_sub571\;
                end if;
              when others =>
                
              end case;
            when pause_getII2227 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v177\ := \$arr1869_value\;
              \$v2224\ := \$v177\;
              \$v2225\ := \$v2224\(0 to 3);
              \$v2219\ := \$v2224\(4 to 67);
              case \$v2225\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2218\ := \$arr1869_ptr_take\;
                if \$v2218\(0) = '1' then
                  state_var2549 <= q_wait2217;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2215;
                end if;
              when "0011" =>
                \$113_p\ := \$v2219\(0 to 4);
                \$v2221\ := \$113_p\;
                \$v2222\ := \$v2221\(0 to 3);
                \$v2220\ := ""&\$v2221\(4);
                case \$v2222\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2218\ := \$arr1869_ptr_take\;
                if \$v2218\(0) = '1' then
                  state_var2549 <= q_wait2217;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2215;
                end if;
              when "0001" =>
                \$114_n\ := \$v2219\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2218\ := \$arr1869_ptr_take\;
                if \$v2218\(0) = '1' then
                  state_var2549 <= q_wait2217;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2215;
                end if;
              when "0000" =>
                \$115_b\ := \$v2219\(0 to 0);
                \$v2223\ := \$115_b\;
                if \$v2223\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2218\ := \$arr1869_ptr_take\;
                  if \$v2218\(0) = '1' then
                    state_var2549 <= q_wait2217;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2215;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2238 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v174\ := \$arr1869_value\;
              \$v2235\ := \$v174\;
              \$v2236\ := \$v2235\(0 to 3);
              \$v2230\ := \$v2235\(4 to 67);
              case \$v2236\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2229\ := \$arr1869_ptr_take\;
                if \$v2229\(0) = '1' then
                  state_var2549 <= q_wait2228;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2226;
                end if;
              when "0011" =>
                \$113_p\ := \$v2230\(0 to 4);
                \$v2232\ := \$113_p\;
                \$v2233\ := \$v2232\(0 to 3);
                \$v2231\ := ""&\$v2232\(4);
                case \$v2233\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2229\ := \$arr1869_ptr_take\;
                if \$v2229\(0) = '1' then
                  state_var2549 <= q_wait2228;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2226;
                end if;
              when "0001" =>
                \$114_n\ := \$v2230\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2229\ := \$arr1869_ptr_take\;
                if \$v2229\(0) = '1' then
                  state_var2549 <= q_wait2228;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2226;
                end if;
              when "0000" =>
                \$115_b\ := \$v2230\(0 to 0);
                \$v2234\ := \$115_b\;
                if \$v2234\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2229\ := \$arr1869_ptr_take\;
                  if \$v2229\(0) = '1' then
                    state_var2549 <= q_wait2228;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2226;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2245 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v167\ := \$arr1869_value\;
              \$v2242\ := \$v167\;
              \$v2243\ := \$v2242\(0 to 3);
              \$v2241\ := \$v2242\(4 to 67);
              case \$v2243\ is
              when "0001" =>
                a := \$v2241\(0 to 31);
                debut := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2240\ := \$arr1869_ptr_take\;
                if \$v2240\(0) = '1' then
                  state_var2549 <= q_wait2239;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2237;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$120_forever5741859\;
              end case;
            when pause_getII2261 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v219\ := \$arr1869_value\;
              \$v2258\ := \$v219\;
              \$v2259\ := \$v2258\(0 to 3);
              \$v2253\ := \$v2258\(4 to 67);
              case \$v2259\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$148_add572\;
              when "0011" =>
                \$113_p\ := \$v2253\(0 to 4);
                \$v2255\ := \$113_p\;
                \$v2256\ := \$v2255\(0 to 3);
                \$v2254\ := ""&\$v2255\(4);
                case \$v2256\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$148_add572\;
              when "0001" =>
                \$114_n\ := \$v2253\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                state_var2549 <= \$148_add572\;
              when "0000" =>
                \$115_b\ := \$v2253\(0 to 0);
                \$v2257\ := \$115_b\;
                if \$v2257\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add572_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$148_add572\;
                end if;
              when others =>
                
              end case;
            when pause_getII2272 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v212\ := \$arr1869_value\;
              \$v2269\ := \$v212\;
              \$v2270\ := \$v2269\(0 to 3);
              \$v2264\ := \$v2269\(4 to 67);
              case \$v2270\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2263\ := \$arr1869_ptr_take\;
                if \$v2263\(0) = '1' then
                  state_var2549 <= q_wait2262;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2260;
                end if;
              when "0011" =>
                \$113_p\ := \$v2264\(0 to 4);
                \$v2266\ := \$113_p\;
                \$v2267\ := \$v2266\(0 to 3);
                \$v2265\ := ""&\$v2266\(4);
                case \$v2267\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2263\ := \$arr1869_ptr_take\;
                if \$v2263\(0) = '1' then
                  state_var2549 <= q_wait2262;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2260;
                end if;
              when "0001" =>
                \$114_n\ := \$v2264\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2263\ := \$arr1869_ptr_take\;
                if \$v2263\(0) = '1' then
                  state_var2549 <= q_wait2262;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2260;
                end if;
              when "0000" =>
                \$115_b\ := \$v2264\(0 to 0);
                \$v2268\ := \$115_b\;
                if \$v2268\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2263\ := \$arr1869_ptr_take\;
                  if \$v2263\(0) = '1' then
                    state_var2549 <= q_wait2262;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2260;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2283 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v209\ := \$arr1869_value\;
              \$v2280\ := \$v209\;
              \$v2281\ := \$v2280\(0 to 3);
              \$v2275\ := \$v2280\(4 to 67);
              case \$v2281\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2274\ := \$arr1869_ptr_take\;
                if \$v2274\(0) = '1' then
                  state_var2549 <= q_wait2273;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2271;
                end if;
              when "0011" =>
                \$113_p\ := \$v2275\(0 to 4);
                \$v2277\ := \$113_p\;
                \$v2278\ := \$v2277\(0 to 3);
                \$v2276\ := ""&\$v2277\(4);
                case \$v2278\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2274\ := \$arr1869_ptr_take\;
                if \$v2274\(0) = '1' then
                  state_var2549 <= q_wait2273;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2271;
                end if;
              when "0001" =>
                \$114_n\ := \$v2275\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2274\ := \$arr1869_ptr_take\;
                if \$v2274\(0) = '1' then
                  state_var2549 <= q_wait2273;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                  state_var2549 <= pause_getI2271;
                end if;
              when "0000" =>
                \$115_b\ := \$v2275\(0 to 0);
                \$v2279\ := \$115_b\;
                if \$v2279\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2274\ := \$arr1869_ptr_take\;
                  if \$v2274\(0) = '1' then
                    state_var2549 <= q_wait2273;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                    state_var2549 <= pause_getI2271;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2291 =>
              \$arr1869_ptr_take\(0) := '0';
              \value\ := \$arr1869_value\;
              \$v2288\ := \value\;
              \$v2289\ := \$v2288\(0 to 3);
              \$v1968\ := \$v2288\(4 to 67);
              case \$v2289\ is
              when "0100" =>
                \$v1178\ := \$v1968\(0 to 63);
                \$v2047\ := \$arr1868_ptr_take\;
                if \$v2047\(0) = '1' then
                  state_var2549 <= q_wait2046;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$v2043\ := \$149_vm_run_code547_arg\(32 to 63);
                  \$arr1868_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                  \$arr1868_write_request\ <= '1';
                  \$arr1868_write\ <= "0001" & \$v2043\&X"00000000";
                  state_var2549 <= pause_setI2044;
                end if;
              when "0011" =>
                p := \$v1968\(0 to 4);
                \$v2286\ := p;
                \$v2287\ := \$v2286\(0 to 3);
                \$v2048\ := ""&\$v2286\(4);
                case \$v2287\ is
                when "0101" =>
                  \$v2073\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v2073\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2549 <= \$120_forever5741850\;
                  else
                    \$v2072\ := \$arr1869_ptr_take\;
                    if \$v2072\(0) = '1' then
                      state_var2549 <= q_wait2071;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                      state_var2549 <= pause_getI2069;
                    end if;
                  end if;
                when "0110" =>
                  \$v2134\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v2134\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2549 <= \$120_forever5741853\;
                  else
                    \$v2133\ := \$arr1869_ptr_take\;
                    if \$v2133\(0) = '1' then
                      state_var2549 <= q_wait2132;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2549 <= pause_getI2130;
                    end if;
                  end if;
                when "0100" =>
                  \$v2153\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v2153\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2549 <= \$120_forever5741856\;
                  else
                    \$v2152\ := \$arr1869_ptr_take\;
                    if \$v2152\(0) = '1' then
                      state_var2549 <= q_wait2151;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2549 <= pause_getI2149;
                    end if;
                  end if;
                when "0011" =>
                  \$v2165\ := eclat_lt(\$192_n\ & "00000000000000000000000000000001");
                  if \$v2165\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("pas assez d'arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2549 <= \$120_forever5741858\;
                  else
                    \$v2164\ := \$arr1869_ptr_take\;
                    if \$v2164\(0) = '1' then
                      state_var2549 <= q_wait2163;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                      state_var2549 <= pause_getI2161;
                    end if;
                  end if;
                when "0010" =>
                  \$146_mul570_arg\ := \$192_n\ & "00000000000000000000000000000001" & \$149_vm_run_code547_arg\(0 to 31);
                  state_var2549 <= \$146_mul570\;
                when "0001" =>
                  \$v2248\ := eclat_lt(\$192_n\ & "00000000000000000000000000000010");
                  if \$v2248\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut 2 arguments pour la soustraction"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2549 <= \$120_forever5741860\;
                  else
                    \$v2247\ := \$arr1869_ptr_take\;
                    if \$v2247\(0) = '1' then
                      state_var2549 <= q_wait2246;
                    else
                      \$arr1869_ptr_take\(0) := '1';
                      \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                      state_var2549 <= pause_getI2244;
                    end if;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2285\ := \$arr1869_ptr_take\;
                  if \$v2285\(0) = '1' then
                    state_var2549 <= q_wait2284;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2282;
                  end if;
                when others =>
                  \$165\ := \$149_vm_run_code547_arg\(0 to 293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                end case;
              when others =>
                \$165\ := \$149_vm_run_code547_arg\(0 to 293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              end case;
            when pause_getII2304 =>
              \$arr1872_ptr_take\(0) := '0';
              \$v1701\ := \$arr1872_value\;
              \$v2302\ := \$arr1869_ptr_take\;
              if \$v2302\(0) = '1' then
                state_var2549 <= q_wait2301;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$v1701\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= v;
                state_var2549 <= pause_setI2299;
              end if;
            when pause_getII2308 =>
              \$arr1869_ptr_take\(0) := '0';
              v := \$arr1869_value\;
              \$v2306\ := \$arr1872_ptr_take\;
              if \$v2306\(0) = '1' then
                state_var2549 <= q_wait2305;
              else
                \$arr1872_ptr_take\(0) := '1';
                \$arr1872_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                state_var2549 <= pause_getI2303;
              end if;
            when pause_getII2315 =>
              \$arr1869_ptr_take\(0) := '0';
              v := \$arr1869_value\;
              \$v2312\ := v;
              \$v2313\ := \$v2312\(0 to 3);
              \$v2311\ := \$v2312\(4 to 67);
              case \$v2313\ is
              when "0000" =>
                x := \$v2311\(0 to 0);
                condition := x;
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & 
                eclat_if(condition & \$149_vm_run_code547_arg\(64 to 95) & eclat_sub(\$195_l\ & "00000000000000000000000000000001")) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when others =>
                condition := eclat_false;
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & 
                eclat_if(condition & \$149_vm_run_code547_arg\(64 to 95) & eclat_sub(\$195_l\ & "00000000000000000000000000000001")) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              end case;
            when pause_getII2322 =>
              \$arr1869_ptr_take\(0) := '0';
              v := \$arr1869_value\;
              \$v2319\ := v;
              \$v2320\ := \$v2319\(0 to 3);
              \$v2318\ := \$v2319\(4 to 67);
              case \$v2320\ is
              when "0000" =>
                x := \$v2318\(0 to 0);
                cond := x;
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$196_l\ & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95)) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when others =>
                cond := eclat_false;
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$196_l\ & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95)) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              end case;
            when pause_getII2330 =>
              \$arr1869_ptr_take\(0) := '0';
              var := \$arr1869_value\;
              \$v2328\ := \$arr1868_ptr_take\;
              if \$v2328\(0) = '1' then
                state_var2549 <= q_wait2327;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$197_i\)));
                \$arr1868_write_request\ <= '1';
                \$arr1868_write\ <= var;
                state_var2549 <= pause_setI2325;
              end if;
            when pause_getII2338 =>
              \$arr1868_ptr_take\(0) := '0';
              local_value := \$arr1868_value\;
              \$v2336\ := \$arr1869_ptr_take\;
              if \$v2336\(0) = '1' then
                state_var2549 <= q_wait2335;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= local_value;
                state_var2549 <= pause_setI2333;
              end if;
            when pause_getII2349 =>
              \$arr1868_ptr_take\(0) := '0';
              \$v247\ := \$arr1868_value\;
              \$v2346\ := \$v247\;
              \$v2347\ := \$v2346\(0 to 3);
              \$v2341\ := \$v2346\(4 to 67);
              case \$v2347\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2340\ := \$arr1868_ptr_take\;
                if \$v2340\(0) = '1' then
                  state_var2549 <= q_wait2339;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2337;
                end if;
              when "0011" =>
                \$113_p\ := \$v2341\(0 to 4);
                \$v2343\ := \$113_p\;
                \$v2344\ := \$v2343\(0 to 3);
                \$v2342\ := ""&\$v2343\(4);
                case \$v2344\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2340\ := \$arr1868_ptr_take\;
                if \$v2340\(0) = '1' then
                  state_var2549 <= q_wait2339;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2337;
                end if;
              when "0001" =>
                \$114_n\ := \$v2341\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v2340\ := \$arr1868_ptr_take\;
                if \$v2340\(0) = '1' then
                  state_var2549 <= q_wait2339;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2337;
                end if;
              when "0000" =>
                \$115_b\ := \$v2341\(0 to 0);
                \$v2345\ := \$115_b\;
                if \$v2345\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2340\ := \$arr1868_ptr_take\;
                  if \$v2340\(0) = '1' then
                    state_var2549 <= q_wait2339;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2337;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2360 =>
              \$arr1868_ptr_take\(0) := '0';
              \$v244\ := \$arr1868_value\;
              \$v2357\ := \$v244\;
              \$v2358\ := \$v2357\(0 to 3);
              \$v2352\ := \$v2357\(4 to 67);
              case \$v2358\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2351\ := \$arr1868_ptr_take\;
                if \$v2351\(0) = '1' then
                  state_var2549 <= q_wait2350;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2348;
                end if;
              when "0011" =>
                \$113_p\ := \$v2352\(0 to 4);
                \$v2354\ := \$113_p\;
                \$v2355\ := \$v2354\(0 to 3);
                \$v2353\ := ""&\$v2354\(4);
                case \$v2355\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2351\ := \$arr1868_ptr_take\;
                if \$v2351\(0) = '1' then
                  state_var2549 <= q_wait2350;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2348;
                end if;
              when "0001" =>
                \$114_n\ := \$v2352\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2351\ := \$arr1868_ptr_take\;
                if \$v2351\(0) = '1' then
                  state_var2549 <= q_wait2350;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                  state_var2549 <= pause_getI2348;
                end if;
              when "0000" =>
                \$115_b\ := \$v2352\(0 to 0);
                \$v2356\ := \$115_b\;
                if \$v2356\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("Fetch["));
                  
                  eclat_print_int(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2351\ := \$arr1868_ptr_take\;
                  if \$v2351\(0) = '1' then
                    state_var2549 <= q_wait2350;
                  else
                    \$arr1868_ptr_take\(0) := '1';
                    \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                    state_var2549 <= pause_getI2348;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2368 =>
              \$arr1870_ptr_take\(0) := '0';
              \$v251\ := \$arr1870_value\;
              \$v2366\ := \$arr1869_ptr_take\;
              if \$v2366\(0) = '1' then
                state_var2549 <= q_wait2365;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= \$v251\;
                state_var2549 <= pause_setI2363;
              end if;
            when pause_getII2376 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v255\ := \$arr1869_value\;
              \$v2374\ := \$arr1870_ptr_take\;
              if \$v2374\(0) = '1' then
                state_var2549 <= q_wait2373;
              else
                \$arr1870_ptr_take\(0) := '1';
                \$arr1870_ptr_write\ <= to_integer(unsigned(\$201_i\));
                \$arr1870_write_request\ <= '1';
                \$arr1870_write\ <= \$v255\;
                state_var2549 <= pause_setI2371;
              end if;
            when pause_getII2387 =>
              \$arr1869_ptr_take\(0) := '0';
              \$v263\ := \$arr1869_value\;
              \$v2384\ := \$v263\;
              \$v2385\ := \$v2384\(0 to 3);
              \$v2379\ := \$v2384\(4 to 67);
              case \$v2385\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0011" =>
                \$113_p\ := \$v2379\(0 to 4);
                \$v2381\ := \$113_p\;
                \$v2382\ := \$v2381\(0 to 3);
                \$v2380\ := ""&\$v2381\(4);
                case \$v2382\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0001" =>
                \$114_n\ := \$v2379\(0 to 31);
                eclat_print_int(\$114_n\);
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0000" =>
                \$115_b\ := \$v2379\(0 to 0);
                \$v2383\ := \$115_b\;
                if \$v2383\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2398 =>
              \$arr1871_ptr_take\(0) := '0';
              \$191_instr\ := \$arr1871_value\;
              \$v2395\ := \$191_instr\;
              \$v2396\ := \$v2395\(0 to 3);
              \$v1967\ := \$v2395\(4 to 71);
              case \$v2396\ is
              when "1000" =>
                \$192_n\ := \$v1967\(0 to 31);
                \$v2293\ := \$arr1869_ptr_take\;
                if \$v2293\(0) = '1' then
                  state_var2549 <= q_wait2292;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2290;
                end if;
              when "0110" =>
                \$193_l\ := \$v1967\(0 to 31);
                \$v2298\ := \$arr1869_ptr_take\;
                if \$v2298\(0) = '1' then
                  state_var2549 <= q_wait2297;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$v2294\ := \$193_l\ & \$149_vm_run_code547_arg\(32 to 63);
                  \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= "0100" & \$v2294\;
                  state_var2549 <= pause_setI2295;
                end if;
              when "1001" =>
                \$v2310\ := \$arr1869_ptr_take\;
                if \$v2310\(0) = '1' then
                  state_var2549 <= q_wait2309;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2307;
                end if;
              when "1100" =>
                \$195_l\ := \$v1967\(0 to 31);
                \$v2317\ := \$arr1869_ptr_take\;
                if \$v2317\(0) = '1' then
                  state_var2549 <= q_wait2316;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2314;
                end if;
              when "1011" =>
                \$196_l\ := \$v1967\(0 to 31);
                \$v2324\ := \$arr1869_ptr_take\;
                if \$v2324\(0) = '1' then
                  state_var2549 <= q_wait2323;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2321;
                end if;
              when "0011" =>
                \$197_i\ := \$v1967\(0 to 31);
                \$v2332\ := \$arr1869_ptr_take\;
                if \$v2332\(0) = '1' then
                  state_var2549 <= q_wait2331;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2329;
                end if;
              when "1010" =>
                \$198_l\ := \$v1967\(0 to 31);
                \$165\ := \$149_vm_run_code547_arg\(0 to 31) & \$149_vm_run_code547_arg\(32 to 63) & eclat_sub(\$198_l\ & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0100" =>
                \$199_i\ := \$v1967\(0 to 31);
                eclat_print_string(of_string("env "));
                
                eclat_print_int(\$149_vm_run_code547_arg\(32 to 63));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(\$149_vm_run_code547_arg\(32 to 63));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2362\ := \$arr1868_ptr_take\;
                if \$v2362\(0) = '1' then
                  state_var2549 <= q_wait2361;
                else
                  \$arr1868_ptr_take\(0) := '1';
                  \$arr1868_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                  state_var2549 <= pause_getI2359;
                end if;
              when "0010" =>
                \$200_i\ := \$v1967\(0 to 31);
                \$v2370\ := \$arr1870_ptr_take\;
                if \$v2370\(0) = '1' then
                  state_var2549 <= q_wait2369;
                else
                  \$arr1870_ptr_take\(0) := '1';
                  \$arr1870_ptr\ <= to_integer(unsigned(\$200_i\));
                  state_var2549 <= pause_getI2367;
                end if;
              when "0001" =>
                \$201_i\ := \$v1967\(0 to 31);
                \$v2378\ := \$arr1869_ptr_take\;
                if \$v2378\(0) = '1' then
                  state_var2549 <= q_wait2377;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2549 <= pause_getI2375;
                end if;
              when "0000" =>
                \$165\ := \$149_vm_run_code547_arg\(0 to 31) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & eclat_add(\$149_vm_run_code547_arg\(128 to 159) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0111" =>
                \$v2390\ := eclat_eq(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & "00000000000000000000000000000000");
                if \$v2390\(0) = '1' then
                  \$v2389\ := \$arr1869_ptr_take\;
                  if \$v2389\(0) = '1' then
                    state_var2549 <= q_wait2388;
                  else
                    \$arr1869_ptr_take\(0) := '1';
                    \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2549 <= pause_getI2386;
                  end if;
                else
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                end if;
              when "0101" =>
                \$204_v\ := \$v1967\(0 to 67);
                \$v2394\ := \$arr1869_ptr_take\;
                if \$v2394\(0) = '1' then
                  state_var2549 <= q_wait2393;
                else
                  \$arr1869_ptr_take\(0) := '1';
                  \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                  \$arr1869_write_request\ <= '1';
                  \$arr1869_write\ <= \$204_v\;
                  state_var2549 <= pause_setI2391;
                end if;
              when others =>
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2549 <= \$208_forever5731845\;
              end case;
            when pause_setI1923 =>
              \$arr1868_write_request\ <= '0';
              state_var2549 <= pause_setII1924;
            when pause_setI1969 =>
              \$arr1872_write_request\ <= '0';
              state_var2549 <= pause_setII1970;
            when pause_setI1973 =>
              \$arr1872_write_request\ <= '0';
              state_var2549 <= pause_setII1974;
            when pause_setI2044 =>
              \$arr1868_write_request\ <= '0';
              state_var2549 <= pause_setII2045;
            when pause_setI2049 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2050;
            when pause_setI2083 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2084;
            when pause_setI2135 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2136;
            when pause_setI2154 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2155;
            when pause_setI2166 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2167;
            when pause_setI2204 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2205;
            when pause_setI2249 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2250;
            when pause_setI2295 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2296;
            when pause_setI2299 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2300;
            when pause_setI2325 =>
              \$arr1868_write_request\ <= '0';
              state_var2549 <= pause_setII2326;
            when pause_setI2333 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2334;
            when pause_setI2363 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2364;
            when pause_setI2371 =>
              \$arr1870_write_request\ <= '0';
              state_var2549 <= pause_setII2372;
            when pause_setI2391 =>
              \$arr1869_write_request\ <= '0';
              state_var2549 <= pause_setII2392;
            when pause_setII1924 =>
              \$arr1868_ptr_take\(0) := '0';
              \$143_copy_args_to_heap544_arg\ := eclat_sub(\$143_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$143_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$143_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
              state_var2549 <= \$143_copy_args_to_heap544\;
            when pause_setII1970 =>
              \$arr1872_ptr_take\(0) := '0';
              \$165\ := eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(\$v1178\(32 to 63) & "00000000000000000000000000000001") & eclat_sub(\$v1178\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII1974 =>
              \$arr1872_ptr_take\(0) := '0';
              \$v1972\ := \$arr1872_ptr_take\;
              if \$v1972\(0) = '1' then
                state_var2549 <= q_wait1971;
              else
                \$arr1872_ptr_take\(0) := '1';
                \$arr1872_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1872_write_request\ <= '1';
                \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$v1178\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(96 to 127);
                state_var2549 <= pause_setI1969;
              end if;
            when pause_setII2045 =>
              \$arr1868_ptr_take\(0) := '0';
              eclat_print_string(of_string("stack["));
              
              eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
              
              eclat_print_string(of_string("] <-"));
              
              \$v2042\ := \$arr1869_ptr_take\;
              if \$v2042\(0) = '1' then
                state_var2549 <= q_wait2041;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2039;
              end if;
            when pause_setII2050 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2084 =>
              \$arr1869_ptr_take\(0) := '0';
              eclat_print_string(of_string("ICIIIIIIIII"));
              
              \$v2081\ := eclat_gt(fst_operand & scd_operand);
              \$v2079\ := "0000" & \$v2081\&"000"& X"000000000000000";
              \$v2080\ := \$v2079\(0 to 3);
              \$v2074\ := \$v2079\(4 to 67);
              case \$v2080\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0011" =>
                \$113_p\ := \$v2074\(0 to 4);
                \$v2076\ := \$113_p\;
                \$v2077\ := \$v2076\(0 to 3);
                \$v2075\ := ""&\$v2076\(4);
                case \$v2077\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0001" =>
                \$114_n\ := \$v2074\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                \$v1966\ := ""&\$165\(293);
                if \$v1966\(0) = '1' then
                  \$149_vm_run_code547_result\ := eclat_unit;
                  result1920 := \$149_vm_run_code547_result\;
                  rdy1921 := eclat_true;
                  state_var2549 <= compute1922;
                else
                  \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                  state_var2549 <= \$149_vm_run_code547\;
                end if;
              when "0000" =>
                \$115_b\ := \$v2074\(0 to 0);
                \$v2078\ := \$115_b\;
                if \$v2078\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
                  \$v1966\ := ""&\$165\(293);
                  if \$v1966\(0) = '1' then
                    \$149_vm_run_code547_result\ := eclat_unit;
                    result1920 := \$149_vm_run_code547_result\;
                    rdy1921 := eclat_true;
                    state_var2549 <= compute1922;
                  else
                    \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                    state_var2549 <= \$149_vm_run_code547\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_setII2136 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2155 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2167 =>
              \$arr1869_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2205 =>
              \$arr1869_ptr_take\(0) := '0';
              eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2250 =>
              \$arr1869_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2296 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2300 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$v1701\(0 to 31) & "00000000000000000000000000000001") & \$v1701\(32 to 63) & \$v1701\(64 to 95) & \$v1701\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2326 =>
              \$arr1868_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2334 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2364 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2372 =>
              \$arr1870_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when pause_setII2392 =>
              \$arr1869_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(32 to 63) & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127) & \$149_vm_run_code547_arg\(128 to 159) & \$149_vm_run_code547_arg\(160 to 191) & \$149_vm_run_code547_arg\(192 to 292) & ""&\$149_vm_run_code547_arg\(293);
              \$v1966\ := ""&\$165\(293);
              if \$v1966\(0) = '1' then
                \$149_vm_run_code547_result\ := eclat_unit;
                result1920 := \$149_vm_run_code547_result\;
                rdy1921 := eclat_true;
                state_var2549 <= compute1922;
              else
                \$149_vm_run_code547_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code547_arg\(294);
                state_var2549 <= \$149_vm_run_code547\;
              end if;
            when q_wait1925 =>
              \$v1926\ := \$arr1868_ptr_take\;
              if \$v1926\(0) = '1' then
                state_var2549 <= q_wait1925;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr_write\ <= to_integer(unsigned(\$143_copy_args_to_heap544_arg\(64 to 95)));
                \$arr1868_write_request\ <= '1';
                \$arr1868_write\ <= \$389\;
                state_var2549 <= pause_setI1923;
              end if;
            when q_wait1929 =>
              \$v1930\ := \$arr1869_ptr_take\;
              if \$v1930\(0) = '1' then
                state_var2549 <= q_wait1929;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$143_copy_args_to_heap544_arg\(32 to 63) & \$143_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI1927;
              end if;
            when q_wait1939 =>
              \$v1940\ := \$arr1869_ptr_take\;
              if \$v1940\(0) = '1' then
                state_var2549 <= q_wait1939;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$145_div569_arg\(64 to 95) & "00000000000000000000000000000001") & \$145_div569_arg\(0 to 31))));
                state_var2549 <= pause_getI1937;
              end if;
            when q_wait1947 =>
              \$v1948\ := \$arr1869_ptr_take\;
              if \$v1948\(0) = '1' then
                state_var2549 <= q_wait1947;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_mul570_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_mul570_arg\(0 to 31))));
                state_var2549 <= pause_getI1945;
              end if;
            when q_wait1955 =>
              \$v1956\ := \$arr1869_ptr_take\;
              if \$v1956\(0) = '1' then
                state_var2549 <= q_wait1955;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_sub571_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_sub571_arg\(0 to 31))));
                state_var2549 <= pause_getI1953;
              end if;
            when q_wait1963 =>
              \$v1964\ := \$arr1869_ptr_take\;
              if \$v1964\(0) = '1' then
                state_var2549 <= q_wait1963;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_add572_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_add572_arg\(0 to 31))));
                state_var2549 <= pause_getI1961;
              end if;
            when q_wait1971 =>
              \$v1972\ := \$arr1872_ptr_take\;
              if \$v1972\(0) = '1' then
                state_var2549 <= q_wait1971;
              else
                \$arr1872_ptr_take\(0) := '1';
                \$arr1872_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1872_write_request\ <= '1';
                \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$v1178\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(96 to 127);
                state_var2549 <= pause_setI1969;
              end if;
            when q_wait1975 =>
              \$v1976\ := \$arr1872_ptr_take\;
              if \$v1976\(0) = '1' then
                state_var2549 <= q_wait1975;
              else
                \$arr1872_ptr_take\(0) := '1';
                \$arr1872_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                \$arr1872_write_request\ <= '1';
                \$arr1872_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001") & \$149_vm_run_code547_arg\(64 to 95) & \$149_vm_run_code547_arg\(96 to 127);
                state_var2549 <= pause_setI1973;
              end if;
            when q_wait1986 =>
              \$v1987\ := \$arr1868_ptr_take\;
              if \$v1987\(0) = '1' then
                state_var2549 <= q_wait1986;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000010")));
                state_var2549 <= pause_getI1984;
              end if;
            when q_wait1997 =>
              \$v1998\ := \$arr1868_ptr_take\;
              if \$v1998\(0) = '1' then
                state_var2549 <= q_wait1997;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI1995;
              end if;
            when q_wait2008 =>
              \$v2009\ := \$arr1868_ptr_take\;
              if \$v2009\(0) = '1' then
                state_var2549 <= q_wait2008;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                state_var2549 <= pause_getI2006;
              end if;
            when q_wait2019 =>
              \$v2020\ := \$arr1869_ptr_take\;
              if \$v2020\(0) = '1' then
                state_var2549 <= q_wait2019;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2017;
              end if;
            when q_wait2030 =>
              \$v2031\ := \$arr1869_ptr_take\;
              if \$v2031\(0) = '1' then
                state_var2549 <= q_wait2030;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                state_var2549 <= pause_getI2028;
              end if;
            when q_wait2041 =>
              \$v2042\ := \$arr1869_ptr_take\;
              if \$v2042\(0) = '1' then
                state_var2549 <= q_wait2041;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2039;
              end if;
            when q_wait2046 =>
              \$v2047\ := \$arr1868_ptr_take\;
              if \$v2047\(0) = '1' then
                state_var2549 <= q_wait2046;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$v2043\ := \$149_vm_run_code547_arg\(32 to 63);
                \$arr1868_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                \$arr1868_write_request\ <= '1';
                \$arr1868_write\ <= "0001" & \$v2043\&X"00000000";
                state_var2549 <= pause_setI2044;
              end if;
            when q_wait2051 =>
              \$v2052\ := \$arr1869_ptr_take\;
              if \$v2052\(0) = '1' then
                state_var2549 <= q_wait2051;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0000" & res&"000"& X"000000000000000";
                state_var2549 <= pause_setI2049;
              end if;
            when q_wait2067 =>
              \$v2068\ := \$arr1869_ptr_take\;
              if \$v2068\(0) = '1' then
                state_var2549 <= q_wait2067;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2549 <= pause_getI2065;
              end if;
            when q_wait2071 =>
              \$v2072\ := \$arr1869_ptr_take\;
              if \$v2072\(0) = '1' then
                state_var2549 <= q_wait2071;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2549 <= pause_getI2069;
              end if;
            when q_wait2085 =>
              \$v2086\ := \$arr1869_ptr_take\;
              if \$v2086\(0) = '1' then
                state_var2549 <= q_wait2085;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$v2082\ := eclat_gt(fst_operand & scd_operand);
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0000" & \$v2082\&"000"& X"000000000000000";
                state_var2549 <= pause_setI2083;
              end if;
            when q_wait2096 =>
              \$v2097\ := \$arr1869_ptr_take\;
              if \$v2097\(0) = '1' then
                state_var2549 <= q_wait2096;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2094;
              end if;
            when q_wait2107 =>
              \$v2108\ := \$arr1869_ptr_take\;
              if \$v2108\(0) = '1' then
                state_var2549 <= q_wait2107;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2549 <= pause_getI2105;
              end if;
            when q_wait2118 =>
              \$v2119\ := \$arr1869_ptr_take\;
              if \$v2119\(0) = '1' then
                state_var2549 <= q_wait2118;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2549 <= pause_getI2116;
              end if;
            when q_wait2125 =>
              \$v2126\ := \$arr1869_ptr_take\;
              if \$v2126\(0) = '1' then
                state_var2549 <= q_wait2125;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2549 <= pause_getI2123;
              end if;
            when q_wait2132 =>
              \$v2133\ := \$arr1869_ptr_take\;
              if \$v2133\(0) = '1' then
                state_var2549 <= q_wait2132;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2549 <= pause_getI2130;
              end if;
            when q_wait2137 =>
              \$v2138\ := \$arr1869_ptr_take\;
              if \$v2138\(0) = '1' then
                state_var2549 <= q_wait2137;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0001" & resultat&X"00000000";
                state_var2549 <= pause_setI2135;
              end if;
            when q_wait2144 =>
              \$v2145\ := \$arr1869_ptr_take\;
              if \$v2145\(0) = '1' then
                state_var2549 <= q_wait2144;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2549 <= pause_getI2142;
              end if;
            when q_wait2151 =>
              \$v2152\ := \$arr1869_ptr_take\;
              if \$v2152\(0) = '1' then
                state_var2549 <= q_wait2151;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2549 <= pause_getI2149;
              end if;
            when q_wait2156 =>
              \$v2157\ := \$arr1869_ptr_take\;
              if \$v2157\(0) = '1' then
                state_var2549 <= q_wait2156;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0001" & resultat&X"00000000";
                state_var2549 <= pause_setI2154;
              end if;
            when q_wait2163 =>
              \$v2164\ := \$arr1869_ptr_take\;
              if \$v2164\(0) = '1' then
                state_var2549 <= q_wait2163;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2161;
              end if;
            when q_wait2168 =>
              \$v2169\ := \$arr1869_ptr_take\;
              if \$v2169\(0) = '1' then
                state_var2549 <= q_wait2168;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0001" & resultat&X"00000000";
                state_var2549 <= pause_setI2166;
              end if;
            when q_wait2179 =>
              \$v2180\ := \$arr1869_ptr_take\;
              if \$v2180\(0) = '1' then
                state_var2549 <= q_wait2179;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2177;
              end if;
            when q_wait2190 =>
              \$v2191\ := \$arr1869_ptr_take\;
              if \$v2191\(0) = '1' then
                state_var2549 <= q_wait2190;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                state_var2549 <= pause_getI2188;
              end if;
            when q_wait2201 =>
              \$v2202\ := \$arr1869_ptr_take\;
              if \$v2202\(0) = '1' then
                state_var2549 <= q_wait2201;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2199;
              end if;
            when q_wait2206 =>
              \$v2207\ := \$arr1869_ptr_take\;
              if \$v2207\(0) = '1' then
                state_var2549 <= q_wait2206;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$v2203\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0001" & \$v2203\&X"00000000";
                state_var2549 <= pause_setI2204;
              end if;
            when q_wait2217 =>
              \$v2218\ := \$arr1869_ptr_take\;
              if \$v2218\(0) = '1' then
                state_var2549 <= q_wait2217;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2215;
              end if;
            when q_wait2228 =>
              \$v2229\ := \$arr1869_ptr_take\;
              if \$v2229\(0) = '1' then
                state_var2549 <= q_wait2228;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                state_var2549 <= pause_getI2226;
              end if;
            when q_wait2239 =>
              \$v2240\ := \$arr1869_ptr_take\;
              if \$v2240\(0) = '1' then
                state_var2549 <= q_wait2239;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2237;
              end if;
            when q_wait2246 =>
              \$v2247\ := \$arr1869_ptr_take\;
              if \$v2247\(0) = '1' then
                state_var2549 <= q_wait2246;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2244;
              end if;
            when q_wait2251 =>
              \$v2252\ := \$arr1869_ptr_take\;
              if \$v2252\(0) = '1' then
                state_var2549 <= q_wait2251;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0001" & resultat&X"00000000";
                state_var2549 <= pause_setI2249;
              end if;
            when q_wait2262 =>
              \$v2263\ := \$arr1869_ptr_take\;
              if \$v2263\(0) = '1' then
                state_var2549 <= q_wait2262;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2260;
              end if;
            when q_wait2273 =>
              \$v2274\ := \$arr1869_ptr_take\;
              if \$v2274\(0) = '1' then
                state_var2549 <= q_wait2273;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\)));
                state_var2549 <= pause_getI2271;
              end if;
            when q_wait2284 =>
              \$v2285\ := \$arr1869_ptr_take\;
              if \$v2285\(0) = '1' then
                state_var2549 <= q_wait2284;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2282;
              end if;
            when q_wait2292 =>
              \$v2293\ := \$arr1869_ptr_take\;
              if \$v2293\(0) = '1' then
                state_var2549 <= q_wait2292;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2290;
              end if;
            when q_wait2297 =>
              \$v2298\ := \$arr1869_ptr_take\;
              if \$v2298\(0) = '1' then
                state_var2549 <= q_wait2297;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$v2294\ := \$193_l\ & \$149_vm_run_code547_arg\(32 to 63);
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= "0100" & \$v2294\;
                state_var2549 <= pause_setI2295;
              end if;
            when q_wait2301 =>
              \$v2302\ := \$arr1869_ptr_take\;
              if \$v2302\(0) = '1' then
                state_var2549 <= q_wait2301;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$v1701\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= v;
                state_var2549 <= pause_setI2299;
              end if;
            when q_wait2305 =>
              \$v2306\ := \$arr1872_ptr_take\;
              if \$v2306\(0) = '1' then
                state_var2549 <= q_wait2305;
              else
                \$arr1872_ptr_take\(0) := '1';
                \$arr1872_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(96 to 127)));
                state_var2549 <= pause_getI2303;
              end if;
            when q_wait2309 =>
              \$v2310\ := \$arr1869_ptr_take\;
              if \$v2310\(0) = '1' then
                state_var2549 <= q_wait2309;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2307;
              end if;
            when q_wait2316 =>
              \$v2317\ := \$arr1869_ptr_take\;
              if \$v2317\(0) = '1' then
                state_var2549 <= q_wait2316;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2314;
              end if;
            when q_wait2323 =>
              \$v2324\ := \$arr1869_ptr_take\;
              if \$v2324\(0) = '1' then
                state_var2549 <= q_wait2323;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2321;
              end if;
            when q_wait2327 =>
              \$v2328\ := \$arr1868_ptr_take\;
              if \$v2328\(0) = '1' then
                state_var2549 <= q_wait2327;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$197_i\)));
                \$arr1868_write_request\ <= '1';
                \$arr1868_write\ <= var;
                state_var2549 <= pause_setI2325;
              end if;
            when q_wait2331 =>
              \$v2332\ := \$arr1869_ptr_take\;
              if \$v2332\(0) = '1' then
                state_var2549 <= q_wait2331;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2329;
              end if;
            when q_wait2335 =>
              \$v2336\ := \$arr1869_ptr_take\;
              if \$v2336\(0) = '1' then
                state_var2549 <= q_wait2335;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= local_value;
                state_var2549 <= pause_setI2333;
              end if;
            when q_wait2339 =>
              \$v2340\ := \$arr1868_ptr_take\;
              if \$v2340\(0) = '1' then
                state_var2549 <= q_wait2339;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                state_var2549 <= pause_getI2337;
              end if;
            when q_wait2350 =>
              \$v2351\ := \$arr1868_ptr_take\;
              if \$v2351\(0) = '1' then
                state_var2549 <= q_wait2350;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code547_arg\(32 to 63) & \$199_i\)));
                state_var2549 <= pause_getI2348;
              end if;
            when q_wait2361 =>
              \$v2362\ := \$arr1868_ptr_take\;
              if \$v2362\(0) = '1' then
                state_var2549 <= q_wait2361;
              else
                \$arr1868_ptr_take\(0) := '1';
                \$arr1868_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(32 to 63)));
                state_var2549 <= pause_getI2359;
              end if;
            when q_wait2365 =>
              \$v2366\ := \$arr1869_ptr_take\;
              if \$v2366\(0) = '1' then
                state_var2549 <= q_wait2365;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= \$v251\;
                state_var2549 <= pause_setI2363;
              end if;
            when q_wait2369 =>
              \$v2370\ := \$arr1870_ptr_take\;
              if \$v2370\(0) = '1' then
                state_var2549 <= q_wait2369;
              else
                \$arr1870_ptr_take\(0) := '1';
                \$arr1870_ptr\ <= to_integer(unsigned(\$200_i\));
                state_var2549 <= pause_getI2367;
              end if;
            when q_wait2373 =>
              \$v2374\ := \$arr1870_ptr_take\;
              if \$v2374\(0) = '1' then
                state_var2549 <= q_wait2373;
              else
                \$arr1870_ptr_take\(0) := '1';
                \$arr1870_ptr_write\ <= to_integer(unsigned(\$201_i\));
                \$arr1870_write_request\ <= '1';
                \$arr1870_write\ <= \$v255\;
                state_var2549 <= pause_setI2371;
              end if;
            when q_wait2377 =>
              \$v2378\ := \$arr1869_ptr_take\;
              if \$v2378\(0) = '1' then
                state_var2549 <= q_wait2377;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2375;
              end if;
            when q_wait2388 =>
              \$v2389\ := \$arr1869_ptr_take\;
              if \$v2389\(0) = '1' then
                state_var2549 <= q_wait2388;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2549 <= pause_getI2386;
              end if;
            when q_wait2393 =>
              \$v2394\ := \$arr1869_ptr_take\;
              if \$v2394\(0) = '1' then
                state_var2549 <= q_wait2393;
              else
                \$arr1869_ptr_take\(0) := '1';
                \$arr1869_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(0 to 31)));
                \$arr1869_write_request\ <= '1';
                \$arr1869_write\ <= \$204_v\;
                state_var2549 <= pause_setI2391;
              end if;
            when q_wait2399 =>
              \$v2400\ := \$arr1871_ptr_take\;
              if \$v2400\(0) = '1' then
                state_var2549 <= q_wait2399;
              else
                \$arr1871_ptr_take\(0) := '1';
                \$arr1871_ptr\ <= to_integer(unsigned(\$149_vm_run_code547_arg\(64 to 95)));
                state_var2549 <= pause_getI2397;
              end if;
            when compute1922 =>
              rdy1921 := eclat_false;
              eclat_print_string(of_string("START (cy="));
              
              eclat_print_int(\$135_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              \$v2402\ := eclat_unit;
              \$149_vm_run_code547_arg\ := "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & eclat_false & "00000000000000000000000000000000" & "0010" & \$v2402\&"000"& X"000000000000000" & eclat_false & argument;
              state_var2549 <= \$149_vm_run_code547\;
            end case;
            \$v2404\ := eclat_not(rdy1921);
            if \$v2404\(0) = '1' then
              result1920 := eclat_unit;
            end if;
            \$136\ := result1920 & rdy1921;
            \$v1919\ := ""&\$136\(1);
            if \$v1919\(0) = '1' then
              eclat_print_string(of_string("END (cy="));
              
              eclat_print_int(\$135_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              result1873 := eclat_unit;
              eclat_print_newline(eclat_unit);
              
              rdy1874 := eclat_true;
              \state\ <= compute1875;
            else
              result1873 := eclat_unit;
              rdy1874 := eclat_true;
              \state\ <= compute1875;
            end if;
          end case;
          
          result <= result1873;
          rdy <= rdy1874;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
