-- code generated from the following source code:
--   ../vm/fail.ecl
--   ../vm/value.ecl
--   ../vm/ram.ecl
--   ../vm/frames.ecl
--   ../vm/vm.ecl
--   ../vm/main.ecl
--
-- with the following command:
--
--    ./eclat -arg=true -relax -notyB ../vm/fail.ecl ../vm/value.ecl ../vm/ram.ecl ../vm/frames.ecl ../vm/vm.ecl ../vm/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute1650, \$128_copy_args_to_heap544\, \$129_pow569\, \$130_div570\, \$131_mul571\, \$132_sub572\, \$133_add573\, \$644_forever5751612\, \$669_forever5751611\, \$694_forever5751610\, \$718_forever5751608\, \$727_forever5751609\, pause_getI1658, pause_getI1666, pause_getI1676, pause_getI1684, pause_getI1692, pause_getI1700, pause_getII1659, pause_getII1667, pause_getII1677, pause_getII1685, pause_getII1693, pause_getII1701, pause_setI1662, pause_setII1663, q_wait1660, q_wait1664, q_wait1668, q_wait1678, q_wait1686, q_wait1694, q_wait1702);
  signal \state\: t_state;
  type t_state_var2261 is (compute2113, \$415_copy_args_to_heap544\, \$416_pow569\, \$417_div570\, \$418_mul571\, \$419_sub572\, \$420_add573\, \$477_forever5751642\, \$481_forever5751636\, \$506_forever5751641\, \$510_forever5751636\, \$535_forever5751640\, \$539_forever5751636\, \$563_forever5751638\, \$567_forever5751636\, \$576_forever5751639\, \$580_forever5751636\, pause_getI2121, pause_getI2129, pause_getI2139, pause_getI2147, pause_getI2155, pause_getI2163, pause_getII2122, pause_getII2130, pause_getII2140, pause_getII2148, pause_getII2156, pause_getII2164, pause_setI2125, pause_setI2169, pause_setI2174, pause_setI2179, pause_setI2185, pause_setI2191, pause_setI2196, pause_setI2201, pause_setI2206, pause_setI2212, pause_setI2217, pause_setI2222, pause_setI2229, pause_setI2234, pause_setI2239, pause_setI2244, pause_setI2249, pause_setII2126, pause_setII2170, pause_setII2175, pause_setII2180, pause_setII2186, pause_setII2192, pause_setII2197, pause_setII2202, pause_setII2207, pause_setII2213, pause_setII2218, pause_setII2223, pause_setII2230, pause_setII2235, pause_setII2240, pause_setII2245, pause_setII2250, q_wait2123, q_wait2127, q_wait2131, q_wait2141, q_wait2149, q_wait2157, q_wait2165, q_wait2171, q_wait2176, q_wait2181, q_wait2187, q_wait2193, q_wait2198, q_wait2203, q_wait2208, q_wait2214, q_wait2219, q_wait2224, q_wait2231, q_wait2236, q_wait2241, q_wait2246, q_wait2251);
  signal state_var2261: t_state_var2261;
  type t_state_var2260 is (compute2110);
  signal state_var2260: t_state_var2260;
  type t_state_var2259 is (compute2105);
  signal state_var2259: t_state_var2259;
  type t_state_var2258 is (compute1708, \$118_forever5741614\, \$118_forever5741621\, \$118_forever5741622\, \$118_forever5741623\, \$118_forever5741624\, \$121_forever5751613\, \$121_forever5751625\, \$121_forever5751626\, \$121_forever5751627\, \$121_forever5751628\, \$121_forever5751629\, \$121_forever5751630\, \$121_forever5751631\, \$121_forever5751632\, \$121_forever5751633\, \$121_forever5751634\, \$121_forever5751635\, \$144_copy_args_to_heap544\, \$145_pow569\, \$146_div570\, \$147_mul571\, \$148_sub572\, \$149_add573\, \$150_vm_run_code547\, \$209_forever5741620\, \$213_forever5741614\, \$259_forever5751619\, \$263_forever5751613\, \$288_forever5751618\, \$292_forever5751613\, \$317_forever5751617\, \$321_forever5751613\, \$345_forever5751615\, \$349_forever5751613\, \$358_forever5751616\, \$362_forever5751613\, pause_getI1716, pause_getI1724, pause_getI1734, pause_getI1742, pause_getI1750, pause_getI1758, pause_getI1796, pause_getI1800, pause_getI1825, pause_getI1836, pause_getI1847, pause_getI1854, pause_getI1861, pause_getI1873, pause_getI1880, pause_getI1892, pause_getI1908, pause_getI1919, pause_getI1930, pause_getI1941, pause_getI1957, pause_getI1968, pause_getI1979, pause_getI1986, pause_getI1999, pause_getI2012, pause_getI2016, pause_getI2023, pause_getI2030, pause_getI2038, pause_getI2046, pause_getI2057, pause_getI2065, pause_getI2073, pause_getI2084, pause_getI2095, pause_getII1717, pause_getII1725, pause_getII1735, pause_getII1743, pause_getII1751, pause_getII1759, pause_getII1797, pause_getII1801, pause_getII1826, pause_getII1837, pause_getII1848, pause_getII1855, pause_getII1862, pause_getII1874, pause_getII1881, pause_getII1893, pause_getII1909, pause_getII1920, pause_getII1931, pause_getII1942, pause_getII1958, pause_getII1969, pause_getII1980, pause_getII1987, pause_getII2000, pause_getII2013, pause_getII2017, pause_getII2024, pause_getII2031, pause_getII2039, pause_getII2047, pause_getII2058, pause_getII2066, pause_getII2074, pause_getII2085, pause_getII2096, pause_setI1720, pause_setI1766, pause_setI1770, pause_setI1775, pause_setI1780, pause_setI1814, pause_setI1866, pause_setI1885, pause_setI1897, pause_setI1946, pause_setI1991, pause_setI2004, pause_setI2008, pause_setI2034, pause_setI2042, pause_setI2061, pause_setI2069, pause_setI2089, pause_setII1721, pause_setII1767, pause_setII1771, pause_setII1776, pause_setII1781, pause_setII1815, pause_setII1867, pause_setII1886, pause_setII1898, pause_setII1947, pause_setII1992, pause_setII2005, pause_setII2009, pause_setII2035, pause_setII2043, pause_setII2062, pause_setII2070, pause_setII2090, q_wait1718, q_wait1722, q_wait1726, q_wait1736, q_wait1744, q_wait1752, q_wait1760, q_wait1768, q_wait1772, q_wait1777, q_wait1782, q_wait1798, q_wait1802, q_wait1816, q_wait1827, q_wait1838, q_wait1849, q_wait1856, q_wait1863, q_wait1868, q_wait1875, q_wait1882, q_wait1887, q_wait1894, q_wait1899, q_wait1910, q_wait1921, q_wait1932, q_wait1943, q_wait1948, q_wait1959, q_wait1970, q_wait1981, q_wait1988, q_wait1993, q_wait2001, q_wait2006, q_wait2010, q_wait2014, q_wait2018, q_wait2025, q_wait2032, q_wait2036, q_wait2040, q_wait2044, q_wait2048, q_wait2059, q_wait2063, q_wait2067, q_wait2071, q_wait2075, q_wait2086, q_wait2091, q_wait2097);
  signal state_var2258: t_state_var2258;
  type array_value_68 is array (natural range <>) of value(0 to 67);
  type array_value_72 is array (natural range <>) of value(0 to 71);
  type array_value_128 is array (natural range <>) of value(0 to 127);
  signal arr1643 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1643_value\ : value(0 to 67);
  signal \$arr1643_ptr\ : natural range 0 to 99;
  signal \$arr1643_ptr_write\ : natural range 0 to 99;
  signal \$arr1643_write\ : value(0 to 67);
  signal \$arr1643_write_request\ : std_logic := '0';
  signal arr1644 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1644_value\ : value(0 to 67);
  signal \$arr1644_ptr\ : natural range 0 to 99;
  signal \$arr1644_ptr_write\ : natural range 0 to 99;
  signal \$arr1644_write\ : value(0 to 67);
  signal \$arr1644_write_request\ : std_logic := '0';
  signal arr1645 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1645_value\ : value(0 to 67);
  signal \$arr1645_ptr\ : natural range 0 to 99;
  signal \$arr1645_ptr_write\ : natural range 0 to 99;
  signal \$arr1645_write\ : value(0 to 67);
  signal \$arr1645_write_request\ : std_logic := '0';
  signal arr1646 : array_value_72(0 to 99) := (others => (others => '0'));
  signal \$arr1646_value\ : value(0 to 71);
  signal \$arr1646_ptr\ : natural range 0 to 99;
  signal \$arr1646_ptr_write\ : natural range 0 to 99;
  signal \$arr1646_write\ : value(0 to 71);
  signal \$arr1646_write_request\ : std_logic := '0';
  signal arr1647 : array_value_128(0 to 99) := (others => (others => '0'));
  signal \$arr1647_value\ : value(0 to 127);
  signal \$arr1647_ptr\ : natural range 0 to 99;
  signal \$arr1647_ptr_write\ : natural range 0 to 99;
  signal \$arr1647_write\ : value(0 to 127);
  signal \$arr1647_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1643_write_request\ = '1' then
                    arr1643(\$arr1643_ptr_write\) <= \$arr1643_write\;
                  else
                   \$arr1643_value\ <= arr1643(\$arr1643_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1644_write_request\ = '1' then
                    arr1644(\$arr1644_ptr_write\) <= \$arr1644_write\;
                  else
                   \$arr1644_value\ <= arr1644(\$arr1644_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1645_write_request\ = '1' then
                    arr1645(\$arr1645_ptr_write\) <= \$arr1645_write\;
                  else
                   \$arr1645_value\ <= arr1645(\$arr1645_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1646_write_request\ = '1' then
                    arr1646(\$arr1646_ptr_write\) <= \$arr1646_write\;
                  else
                   \$arr1646_value\ <= arr1646(\$arr1646_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1647_write_request\ = '1' then
                    arr1647(\$arr1647_ptr_write\) <= \$arr1647_write\;
                  else
                   \$arr1647_value\ <= arr1647(\$arr1647_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$137\, \$412\ : value(0 to 1) := (others => '0');
      variable \$147_mul571_arg\, \$148_sub572_arg\, \$132_sub572_arg\, 
               \$128_copy_args_to_heap544_arg\, \$146_div570_arg\, 
               \$144_copy_args_to_heap544_arg\, \$133_add573_arg\, 
               \$418_mul571_arg\, \$415_copy_args_to_heap544_arg\, 
               \$130_div570_arg\, \$416_pow569_arg\, \$145_pow569_arg\, 
               \$419_sub572_arg\, \$149_add573_arg\, \$417_div570_arg\, 
               \$129_pow569_arg\, \$420_add573_arg\, \$131_mul571_arg\ : value(0 to 95) := (others => '0');
      variable \$v1961\, \$v2136\, \$v1755\, \$v1784\, \$v1818\, \$v2077\, 
               \$v1840\, \$v1731\, \$v1747\, \$v1785\, \$v2050\, \$v1923\, 
               \$v1829\, \$v2160\, \$v1934\, \$v1709\, \$v1681\, \$v1673\, 
               \$v1805\, \$v2152\, \$v1739\, \$v2020\, \$v1791\, \$v1870\, 
               \$v2027\, \$v1972\, \$v1137\, \$v1697\, \$v1765\, \$v1912\, 
               \$v2003\, \$v2144\, \$v1877\, \$v1788\, \$v1689\, \$v1858\, 
               \$v1851\, \$v1983\, \$v1651\, \$v2114\, \$v1901\, \$v1950\, 
               \$v1889\ : value(0 to 63) := (others => '0');
      variable \$v2093\, \$192_instr\ : value(0 to 71) := (others => '0');
      variable \$114_p\, \$762_p\, \$v2052\, \$v2227\, \$v1963\, \$v1842\, 
               \$615_p\, \$v1903\, \$v1914\, \$v1925\, \$v1711\, \$v1995\, 
               \$v2079\, \$397_p\, \$v1831\, \$v1974\, \$v1936\, \$v1952\, 
               \$v1653\, \$v2116\, p, \$v1820\, \$v1807\ : value(0 to 4) := (others => '0');
      variable \$v1996\, \$v2146\, \$v1964\, \$v1998\, \$v1953\, \$v1872\, 
               \$v1918\, \$v2080\, \$v2120\, \$v1879\, \$v1675\, \$v1975\, 
               \$v1808\, \$v1915\, \$v2053\, \$v1940\, \$v1929\, \$v1757\, 
               \$v1967\, \$v1860\, \$v1790\, \$v1835\, \$v2022\, \$v2162\, 
               \$v1699\, \$v2083\, \$v1937\, \$v1978\, \$v1654\, \$v1907\, 
               \$v2094\, \$v1832\, \$v1787\, \$v1733\, \$v1811\, \$v2117\, 
               \$v2154\, \$v1683\, \$v1904\, \$v1956\, \$v1853\, \$v1891\, 
               \$v1795\, \$v2056\, \$v1926\, \$v1985\, \$v1741\, \$v1824\, 
               \$v2138\, \$v1715\, \$v1712\, \$v1657\, \$v1846\, \$v1749\, 
               \$v1821\, \$v1793\, \$v1691\, \$v1843\, \$v2029\ : value(0 to 3) := (others => '0');
      variable \$150_vm_run_code547_arg\ : value(0 to 294) := (others => '0');
      variable \$v1476\ : value(0 to 127) := (others => '0');
      variable \$v1916\, \$v1960\, cond, \$v2037\, \$v1809\, \$v1938\, 
               \$v2210\, \$v1944\, \$v1672\, \$116_b\, \$v1769\, \$v1839\, 
               \$v1924\, \$v2107\, \$v2247\, \$v1989\, \$v2209\, \$v1828\, 
               rdy1649, \$150_vm_run_code547_result\, \$v1779\, condition, 
               \$765_b\, rdy1707, \$v1884\, \$v2252\, rdy2109, \$v1745\, 
               \$v2072\, \$v2135\, \$v2199\, \$v2011\, \$v2100\, \$v1696\, 
               \$v1804\, \$v1954\, \$v2188\, \$v2220\, \$v1669\, 
               \$135_is_loaded\, \$v1799\, x, \$v2098\, \$v2142\, \$v1723\, 
               result2108, \$v2254\, \$v2143\, \$v2168\, \$v1896\, \$v2054\, 
               \$v1951\, \$v1705\, result2111, \$v1911\, \$v1935\, \$99_a1\, 
               \$v1976\, \$v1803\, \$v2133\, \$v2002\, \$v1762\, \$410\, 
               \$v2248\, result1706, \$v2118\, \$v2049\, \$v2216\, \$v1883\, 
               \$v1876\, \$v2099\, \$v1713\, \$v1864\, \$v1857\, \$v2051\, 
               \$v1888\, \$v1665\, \$v2128\, \$v1905\, \$v1737\, \$v2194\, 
               res, \$v1729\, \$v2204\, \$v2167\, \$v1965\, \$v2026\, 
               \$v1704\, \$v2172\, \$v1850\, \$v1990\, \$v2257\, \$v2078\, 
               \$v2102\, \$v2158\, \$v2150\, \$v1773\, \$v1761\, \$400_b\, 
               rdy2112, result1648, \$v1900\, \$v2242\, \$v1679\, \$v2132\, 
               \$v2087\, \$v2159\, \$v2081\, \$v2166\, \$v2045\, b2, 
               \$v1913\, \$v1812\, \$v1830\, \$v2041\, \$v1933\, \$v1730\, 
               \$v1728\, \$v1971\, \$v2068\, \$v1738\, \$v2033\, \$v1688\, 
               \$v1822\, \$v1687\, \$v1841\, \$v1895\, \$v2182\, \$v2124\, 
               \$v1753\, \$v1680\, \$v2151\, \$v2255\, \$v1833\, \$v2225\, 
               \$v1710\, \$v1746\, \$v2115\, \$v1727\, \$v2177\, \$v1703\, 
               \$v1902\, \$v2092\, \$v1962\, \$v1754\, \$v1671\, \$v1869\, 
               \$v1719\, \$v1994\, \$v1819\, \$v1778\, \$v1670\, \$v2060\, 
               \$v2076\, \$v2226\, \$v2015\, \$v2088\, \$618_b\, \$v1695\, 
               \$v2232\, \$v1865\, \$v2215\, \$v1817\, \$v1844\, \$v2007\, 
               \$v2205\, \$v1922\, \$v1949\, \$v2134\, \$v2019\, \$v1783\, 
               \$v1927\, \$v1973\, rdy2104, \$v1655\, \$v1661\, \$v2237\, 
               \$v1813\, \$v1806\, \$v1763\, \$v1982\, \$v2064\, \$v1652\ : value(0 to 0) := (others => '0');
      variable \$617_n\, \$336_divisor\, \$497_int_value\, \$554_divisor\, 
               \$408\, \$148_sub572_result\, fst_operand, \$665_a\, \$531_a\, 
               result2103, scd_operand, \$200_i\, base, debut, 
               \$149_add573_result\, \$723_a\, \$v2238\, \$v2189\, \$640_a\, 
               \$279_int_value\, \$468_int_value\, \$146_div570_result\, 
               \$144_copy_args_to_heap544_result\, \$399_n\, \$313_a\, 
               \$526_int_value\, \$197_l\, \$473_a\, \$v2221\, \$115_n\, 
               \$196_l\, \$198_i\, \$193_n\, \$136_cy\, \$201_i\, \$v2195\, 
               \$685_int_value\, \$635_int_value\, \$709_divisor\, \$284_a\, 
               \$308_int_value\, \$199_l\, \$690_a\, \$v2183\, \$v1945\, 
               \$502_a\, \$v2243\, \$v2233\, \$194_l\, \$255_a\, \$100_a\, 
               exponent, \$v2178\, \$v1774\, \$145_pow569_result\, \$572_a\, 
               resultat, \$v2173\, \$v2200\, \$147_mul571_result\, \$764_n\, 
               \$660_int_value\, b, \$250_int_value\, \$354_a\, \$202_i\, a : value(0 to 31) := (others => '0');
      variable \$166\ : value(0 to 293) := (others => '0');
      variable \$v1764\, \$v1698\, \$v1682\, \$v51\, \$v1939\, \$v1794\, 
               \$v229\, \$760\, \$v1748\, \$v2190\, \$v2028\, \$v217\, 
               \$v1997\, \$249_v\, second_value, \$v46\, \$v69\, \$v1834\, 
               first_value, \$v1789\, \$v1871\, \$v160\, \$v221\, \$684_v\, 
               \$v1823\, \$v2055\, \$v2153\, \$v1928\, \$v1732\, \$v1890\, 
               \$v1792\, \$v1878\, \$571\, \$v1859\, \$v93\, \$205_v\, 
               \$v2161\, \$395\, \$v1845\, \$v2211\, \$v2228\, \$v1810\, 
               \$404\, var, \$v125\, \$v2184\, \$v57\, \$v2137\, \$467_v\, 
               \$v1906\, \$722\, \$v48\, \$v1852\, \$v1674\, \$v2145\, 
               \$v1917\, \$v153\, \$278_v\, \$v1690\, \$769\, \$613\, \$353\, 
               \$v150\, \$v1955\, \value\, \$525_v\, \$v1714\, \$v1756\, 
               \$v1966\, \$v2119\, \$307_v\, \$v67\, \$v2082\, \$v115\, 
               \$622\, \$v118\, \$v54\, \$v1786\, \$496_v\, \$v213\, 
               \$659_v\, \$v1977\, \$634_v\, \$v1740\, local_value, \$v1984\, 
               \$v2021\, \$v143\, v, \$v1656\, \$v176\ : value(0 to 67) := (others => '0');
      variable \$arr1643_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1644_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1645_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1646_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1647_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(a); default_zero(\$202_i\); default_zero(\$v1652\); 
          default_zero(\$v2064\); default_zero(\$v1982\); 
          default_zero(\$131_mul571_arg\); default_zero(\$v2029\); 
          default_zero(\$v176\); default_zero(\$v1763\); 
          default_zero(\$v1806\); default_zero(\$v1889\); 
          default_zero(\$420_add573_arg\); default_zero(\$v1813\); 
          default_zero(\$354_a\); default_zero(\$v1843\); 
          default_zero(\$v1656\); default_zero(\$v2237\); 
          default_zero(\$v1661\); default_zero(\$v1691\); 
          default_zero(\$129_pow569_arg\); default_zero(v); 
          default_zero(\$v1655\); default_zero(rdy2104); 
          default_zero(\$v1950\); default_zero(\$v143\); 
          default_zero(\$250_int_value\); default_zero(\$192_instr\); 
          default_zero(\$v1973\); default_zero(\$v1927\); 
          default_zero(\$v1783\); default_zero(b); 
          default_zero(\$660_int_value\); default_zero(\$v2019\); 
          default_zero(\$v1901\); default_zero(\$v2134\); 
          default_zero(\$v1949\); default_zero(\$417_div570_arg\); 
          default_zero(\$v1793\); default_zero(\$v1922\); 
          default_zero(\$v2021\); default_zero(\$v2205\); 
          default_zero(\$v1984\); default_zero(local_value); 
          default_zero(\$v1821\); default_zero(\$v2007\); 
          default_zero(\$v1844\); default_zero(\$v1817\); 
          default_zero(\$v2215\); default_zero(\$764_n\); 
          default_zero(\$v1740\); default_zero(\$v1865\); 
          default_zero(\$147_mul571_result\); default_zero(\$v1749\); 
          default_zero(\$v2232\); default_zero(\$v2114\); 
          default_zero(\$v1651\); default_zero(\$634_v\); 
          default_zero(\$149_add573_arg\); default_zero(\$v2200\); 
          default_zero(\$v1695\); default_zero(\$618_b\); 
          default_zero(\$v1846\); default_zero(\$v1657\); 
          default_zero(\$v2173\); default_zero(\$v1712\); 
          default_zero(\$v1715\); default_zero(\$v2088\); 
          default_zero(\$v2015\); default_zero(\$v1977\); 
          default_zero(\$v2226\); default_zero(\$659_v\); 
          default_zero(\$v2076\); default_zero(\$v213\); 
          default_zero(\$v2060\); default_zero(\$496_v\); 
          default_zero(\$v1670\); default_zero(\$v1778\); 
          default_zero(\$v1983\); default_zero(\$v1786\); 
          default_zero(\$v54\); default_zero(\$v118\); 
          default_zero(\$v1819\); default_zero(\$v1994\); 
          default_zero(\$v1851\); default_zero(resultat); 
          default_zero(\$572_a\); default_zero(\$622\); 
          default_zero(\$145_pow569_result\); default_zero(\$v115\); 
          default_zero(\$v1858\); default_zero(\$v1719\); 
          default_zero(\$v1869\); default_zero(\$v2138\); 
          default_zero(\$v1824\); default_zero(\$v1671\); 
          default_zero(\$v1741\); default_zero(\$v1985\); 
          default_zero(\$v2082\); default_zero(\$v1754\); 
          default_zero(\$v1689\); default_zero(\$v1774\); 
          default_zero(\$v67\); default_zero(\$v1962\); 
          default_zero(\$v2178\); default_zero(\$419_sub572_arg\); 
          default_zero(\$v2092\); default_zero(\$v1926\); 
          default_zero(\$v1902\); default_zero(\$v1807\); 
          default_zero(\$307_v\); default_zero(\$v1703\); 
          default_zero(\$v2119\); default_zero(\$v1966\); 
          default_zero(\$v2177\); default_zero(\$v1756\); 
          default_zero(\$v1714\); default_zero(\$v2056\); 
          default_zero(\$v1788\); default_zero(\$525_v\); 
          default_zero(\$v1727\); default_zero(\$v1795\); 
          default_zero(\$v1877\); default_zero(\$v2115\); 
          default_zero(\$v1820\); default_zero(exponent); 
          default_zero(\$v1746\); default_zero(\$v1891\); 
          default_zero(\$v1710\); default_zero(\$v1853\); 
          default_zero(\$100_a\); default_zero(\$255_a\); 
          default_zero(\$v2225\); default_zero(p); default_zero(\$v1956\); 
          default_zero(\value\); default_zero(\$194_l\); 
          default_zero(\$v1833\); default_zero(\$v2255\); 
          default_zero(\$v2144\); default_zero(\$v2116\); 
          default_zero(\$v2151\); default_zero(\$v1680\); 
          default_zero(\$v1753\); default_zero(\$v2124\); 
          default_zero(\$v2182\); default_zero(\$v1895\); 
          default_zero(\$v1955\); default_zero(\$v1841\); 
          default_zero(\$v1687\); default_zero(\$v2233\); 
          default_zero(\$v150\); default_zero(\$v1653\); 
          default_zero(\$v1904\); default_zero(\$353\); default_zero(\$412\); 
          default_zero(\$v1822\); default_zero(\$v1683\); 
          default_zero(\$v2243\); default_zero(\$v1688\); 
          default_zero(\$v2033\); default_zero(\$v1738\); 
          default_zero(\$145_pow569_arg\); default_zero(\$502_a\); 
          default_zero(\$v2003\); default_zero(\$v1912\); 
          default_zero(\$v2068\); default_zero(\$613\); 
          default_zero(\$v1971\); default_zero(\$769\); 
          default_zero(\$v1728\); default_zero(\$v1730\); 
          default_zero(\$v1933\); default_zero(\$v1690\); 
          default_zero(\$278_v\); default_zero(\$v1945\); 
          default_zero(\$v1765\); default_zero(\$v2041\); 
          default_zero(\$v1830\); default_zero(\$v2183\); 
          default_zero(\$v1812\); default_zero(\$v153\); 
          default_zero(\$v1913\); default_zero(\$v1952\); default_zero(b2); 
          default_zero(\$v2045\); default_zero(\$v1697\); 
          default_zero(\$v2166\); default_zero(\$690_a\); 
          default_zero(\$199_l\); default_zero(\$v1936\); 
          default_zero(\$v1917\); default_zero(\$v2154\); 
          default_zero(\$v2081\); default_zero(\$v2145\); 
          default_zero(\$v2159\); default_zero(\$416_pow569_arg\); 
          default_zero(\$v1674\); default_zero(\$308_int_value\); 
          default_zero(\$v2117\); default_zero(\$v1974\); 
          default_zero(\$130_div570_arg\); default_zero(\$284_a\); 
          default_zero(\$v2087\); default_zero(\$v1811\); 
          default_zero(\$v2132\); default_zero(\$v1137\); 
          default_zero(\$v1972\); default_zero(\$v1733\); 
          default_zero(\$v1679\); default_zero(\$v2027\); 
          default_zero(\$v2242\); default_zero(\$v1852\); 
          default_zero(\$v48\); default_zero(\$v1900\); default_zero(\$722\); 
          default_zero(\$v1906\); 
          default_zero(\$415_copy_args_to_heap544_arg\); 
          default_zero(result1648); default_zero(\$v1787\); 
          default_zero(rdy2112); default_zero(\$v1832\); 
          default_zero(\$709_divisor\); default_zero(\$v1870\); 
          default_zero(\$v1791\); default_zero(\$635_int_value\); 
          default_zero(\$685_int_value\); default_zero(\$467_v\); 
          default_zero(\$v2137\); default_zero(\$v57\); 
          default_zero(\$400_b\); default_zero(\$v2195\); 
          default_zero(\$v1761\); default_zero(\$v1773\); 
          default_zero(\$v2184\); default_zero(\$v125\); 
          default_zero(\$201_i\); default_zero(\$v2094\); 
          default_zero(\$v2150\); default_zero(\$136_cy\); 
          default_zero(\$v1831\); default_zero(\$193_n\); default_zero(var); 
          default_zero(\$v2158\); default_zero(\$v2020\); 
          default_zero(\$397_p\); default_zero(\$v2102\); 
          default_zero(\$198_i\); default_zero(\$196_l\); 
          default_zero(\$v2078\); default_zero(\$115_n\); 
          default_zero(\$v2257\); default_zero(\$v2221\); 
          default_zero(\$404\); default_zero(\$v1739\); 
          default_zero(\$v1990\); default_zero(\$v1850\); 
          default_zero(\$v2172\); default_zero(\$v1810\); 
          default_zero(\$v2228\); default_zero(\$473_a\); 
          default_zero(\$v2152\); default_zero(\$418_mul571_arg\); 
          default_zero(\$v1704\); default_zero(\$v2026\); 
          default_zero(\$v1965\); default_zero(\$v1907\); 
          default_zero(\$v2167\); default_zero(\$v1805\); 
          default_zero(\$v2211\); default_zero(\$v2204\); 
          default_zero(\$v1845\); default_zero(\$v1654\); 
          default_zero(\$v2079\); default_zero(\$v1729\); 
          default_zero(\$v1978\); default_zero(\$v1937\); default_zero(res); 
          default_zero(\$395\); default_zero(\$v2194\); 
          default_zero(\$v2161\); default_zero(\$v1737\); 
          default_zero(\$v1905\); default_zero(\$166\); 
          default_zero(\$v2128\); default_zero(\$v2083\); 
          default_zero(\$v1699\); default_zero(\$197_l\); 
          default_zero(\$v1995\); default_zero(\$v1665\); 
          default_zero(\$v1888\); default_zero(\$v2051\); 
          default_zero(\$v1857\); default_zero(\$v1864\); 
          default_zero(\$v2162\); default_zero(\$v1713\); 
          default_zero(\$v2099\); default_zero(\$526_int_value\); 
          default_zero(\$v1876\); default_zero(\$v1711\); 
          default_zero(\$205_v\); default_zero(\$v1883\); 
          default_zero(\$v1925\); default_zero(\$v2216\); 
          default_zero(\$v2022\); default_zero(\$v93\); 
          default_zero(\$v1859\); default_zero(\$571\); 
          default_zero(\$v2049\); default_zero(\$v1878\); 
          default_zero(\$313_a\); default_zero(\$v2118\); 
          default_zero(\$v1476\); default_zero(\$v1673\); 
          default_zero(\$v1835\); default_zero(\$v1681\); 
          default_zero(result1706); default_zero(\$v1790\); 
          default_zero(\$v2248\); default_zero(\$410\); 
          default_zero(\$v1792\); default_zero(\$v1890\); 
          default_zero(\$v1860\); default_zero(\$v1732\); 
          default_zero(\$v1967\); default_zero(\$v1914\); 
          default_zero(\$v1762\); default_zero(\$v2002\); 
          default_zero(\$v1709\); default_zero(\$v2133\); 
          default_zero(\$v1803\); default_zero(\$v1976\); 
          default_zero(\$99_a1\); default_zero(\$399_n\); 
          default_zero(\$144_copy_args_to_heap544_result\); 
          default_zero(\$v1935\); default_zero(\$146_div570_result\); 
          default_zero(\$133_add573_arg\); default_zero(\$v1934\); 
          default_zero(\$v1911\); default_zero(\$468_int_value\); 
          default_zero(\$v2160\); default_zero(result2111); 
          default_zero(\$v1928\); default_zero(\$279_int_value\); 
          default_zero(\$640_a\); default_zero(\$v1705\); 
          default_zero(\$v1951\); default_zero(\$v2054\); 
          default_zero(\$v1757\); default_zero(\$v1896\); 
          default_zero(\$v1829\); default_zero(\$v2168\); 
          default_zero(\$v2153\); default_zero(\$v2143\); 
          default_zero(\$v1929\); 
          default_zero(\$144_copy_args_to_heap544_arg\); 
          default_zero(\$v2254\); default_zero(result2108); 
          default_zero(\$v2055\); default_zero(\$v1723\); 
          default_zero(\$v2142\); default_zero(\$v2098\); default_zero(x); 
          default_zero(\$v1799\); default_zero(\$v1940\); 
          default_zero(\$v1823\); default_zero(\$135_is_loaded\); 
          default_zero(\$684_v\); default_zero(\$v1669\); 
          default_zero(\$v2220\); default_zero(\$v2188\); 
          default_zero(\$v1954\); default_zero(\$v2189\); 
          default_zero(\$v2238\); default_zero(\$723_a\); 
          default_zero(\$v2053\); default_zero(\$v1903\); 
          default_zero(\$149_add573_result\); default_zero(\$v221\); 
          default_zero(debut); default_zero(\$v1804\); 
          default_zero(\$v1696\); default_zero(\$v1923\); 
          default_zero(\$146_div570_arg\); default_zero(\$v2100\); 
          default_zero(\$v2011\); default_zero(\$v160\); 
          default_zero(\$v1871\); default_zero(\$v2199\); default_zero(base); 
          default_zero(\$v2135\); default_zero(\$v1915\); 
          default_zero(\$v1789\); default_zero(first_value); 
          default_zero(\$v2050\); default_zero(\$v1834\); 
          default_zero(\$v1808\); default_zero(\$v2072\); 
          default_zero(\$200_i\); default_zero(\$v1785\); 
          default_zero(\$615_p\); default_zero(\$v1745\); 
          default_zero(\$v1747\); default_zero(\$v69\); 
          default_zero(\$128_copy_args_to_heap544_arg\); 
          default_zero(\$v1975\); default_zero(rdy2109); 
          default_zero(\$v46\); default_zero(scd_operand); 
          default_zero(second_value); default_zero(\$137\); 
          default_zero(\$249_v\); default_zero(\$v1997\); 
          default_zero(\$v217\); default_zero(\$v2028\); 
          default_zero(\$v2252\); default_zero(\$v1675\); 
          default_zero(result2103); default_zero(\$v1879\); 
          default_zero(\$v1842\); default_zero(\$132_sub572_arg\); 
          default_zero(\$v1884\); default_zero(\$v1963\); 
          default_zero(\$v2190\); default_zero(\$531_a\); 
          default_zero(\$v1731\); default_zero(\$665_a\); 
          default_zero(\$v2227\); default_zero(\$v1748\); 
          default_zero(rdy1707); default_zero(\$v2120\); 
          default_zero(\$765_b\); default_zero(\$v2080\); 
          default_zero(\$v1918\); default_zero(\$v1840\); 
          default_zero(condition); default_zero(fst_operand); 
          default_zero(\$v2052\); default_zero(\$760\); 
          default_zero(\$148_sub572_result\); default_zero(\$v1779\); 
          default_zero(\$150_vm_run_code547_result\); default_zero(\$v229\); 
          default_zero(\$v1794\); default_zero(rdy1649); 
          default_zero(\$v2093\); default_zero(\$v2077\); 
          default_zero(\$762_p\); default_zero(\$v1872\); 
          default_zero(\$148_sub572_arg\); default_zero(\$v1828\); 
          default_zero(\$v2209\); default_zero(\$v1989\); 
          default_zero(\$408\); default_zero(\$v2247\); 
          default_zero(\$v2107\); default_zero(\$v1939\); 
          default_zero(\$v1924\); default_zero(\$v1839\); 
          default_zero(\$v1769\); default_zero(\$v1953\); 
          default_zero(\$116_b\); default_zero(\$147_mul571_arg\); 
          default_zero(\$v1998\); default_zero(\$v1964\); 
          default_zero(\$v51\); default_zero(\$v1672\); 
          default_zero(\$v1944\); default_zero(\$v2210\); 
          default_zero(\$v1938\); default_zero(\$v1818\); 
          default_zero(\$v1682\); default_zero(\$554_divisor\); 
          default_zero(\$v1784\); default_zero(\$497_int_value\); 
          default_zero(\$114_p\); default_zero(\$v1809\); 
          default_zero(\$336_divisor\); default_zero(\$v2146\); 
          default_zero(\$v2037\); default_zero(cond); 
          default_zero(\$150_vm_run_code547_arg\); default_zero(\$v1960\); 
          default_zero(\$v1698\); default_zero(\$v1764\); 
          default_zero(\$v1916\); default_zero(\$617_n\); 
          default_zero(\$v1755\); default_zero(\$v2136\); 
          default_zero(\$v1996\); default_zero(\$v1961\); 
          rdy <= "1";
          rdy1649 := "0";
          \state\ <= compute1650;
          state_var2261 <= compute2113;
          state_var2260 <= compute2110;
          state_var2259 <= compute2105;
          state_var2258 <= compute1708;
          
        else if run = '1' then
          case \state\ is
          when \$128_copy_args_to_heap544\ =>
            \$v1670\ := eclat_eq(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1670\(0) = '1' then
              \state\ <= \$128_copy_args_to_heap544\;
            else
              \$v1669\ := \$arr1644_ptr_take\;
              if \$v1669\(0) = '1' then
                \state\ <= q_wait1668;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$128_copy_args_to_heap544_arg\(32 to 63) & \$128_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                \state\ <= pause_getI1666;
              end if;
            end if;
          when \$129_pow569\ =>
            \$v1671\ := eclat_eq(\$129_pow569_arg\(32 to 63) & "00000000000000000000000000000000");
            if \$v1671\(0) = '1' then
              \state\ <= \$129_pow569\;
            else
              \$129_pow569_arg\ := \$129_pow569_arg\(0 to 31) & eclat_sub(\$129_pow569_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$129_pow569_arg\(64 to 95) & \$129_pow569_arg\(0 to 31));
              \state\ <= \$129_pow569\;
            end if;
          when \$130_div570\ =>
            \$v1680\ := eclat_eq(\$130_div570_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1680\(0) = '1' then
              \state\ <= \$130_div570\;
            else
              \$v1679\ := \$arr1644_ptr_take\;
              if \$v1679\(0) = '1' then
                \state\ <= q_wait1678;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_div570_arg\(0 to 31))));
                \state\ <= pause_getI1676;
              end if;
            end if;
          when \$131_mul571\ =>
            \$v1688\ := eclat_eq(\$131_mul571_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1688\(0) = '1' then
              \state\ <= \$131_mul571\;
            else
              \$v1687\ := \$arr1644_ptr_take\;
              if \$v1687\(0) = '1' then
                \state\ <= q_wait1686;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_mul571_arg\(0 to 31))));
                \state\ <= pause_getI1684;
              end if;
            end if;
          when \$132_sub572\ =>
            \$v1696\ := eclat_eq(\$132_sub572_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1696\(0) = '1' then
              \state\ <= \$132_sub572\;
            else
              \$v1695\ := \$arr1644_ptr_take\;
              if \$v1695\(0) = '1' then
                \state\ <= q_wait1694;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_sub572_arg\(0 to 31))));
                \state\ <= pause_getI1692;
              end if;
            end if;
          when \$133_add573\ =>
            \$v1704\ := eclat_eq(\$133_add573_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1704\(0) = '1' then
              \state\ <= \$133_add573\;
            else
              \$v1703\ := \$arr1644_ptr_take\;
              if \$v1703\(0) = '1' then
                \state\ <= q_wait1702;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$133_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$133_add573_arg\(0 to 31))));
                \state\ <= pause_getI1700;
              end if;
            end if;
          when \$644_forever5751612\ =>
            \state\ <= \$644_forever5751612\;
          when \$669_forever5751611\ =>
            \state\ <= \$669_forever5751611\;
          when \$694_forever5751610\ =>
            \state\ <= \$694_forever5751610\;
          when \$718_forever5751608\ =>
            \state\ <= \$718_forever5751608\;
          when \$727_forever5751609\ =>
            \state\ <= \$727_forever5751609\;
          when pause_getI1658 =>
            \state\ <= pause_getII1659;
          when pause_getI1666 =>
            \state\ <= pause_getII1667;
          when pause_getI1676 =>
            \state\ <= pause_getII1677;
          when pause_getI1684 =>
            \state\ <= pause_getII1685;
          when pause_getI1692 =>
            \state\ <= pause_getII1693;
          when pause_getI1700 =>
            \state\ <= pause_getII1701;
          when pause_getII1659 =>
            \$arr1644_ptr_take\(0) := '0';
            \$760\ := \$arr1644_value\;
            \$v1656\ := \$760\;
            \$v1657\ := \$v1656\(0 to 3);
            \$v1651\ := \$v1656\(4 to 67);
            case \$v1657\ is
            when "0100" =>
              eclat_print_string(of_string("fermeture"));
              
              eclat_print_newline(eclat_unit);
              
              \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
              \state\ <= \$128_copy_args_to_heap544\;
            when "0011" =>
              \$762_p\ := \$v1651\(0 to 4);
              \$v1653\ := \$762_p\;
              \$v1654\ := \$v1653\(0 to 3);
              \$v1652\ := ""&\$v1653\(4);
              case \$v1654\ is
              when "0110" =>
                eclat_print_string(of_string("<"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0101" =>
                eclat_print_string(of_string("=="));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0100" =>
                eclat_print_string(of_string("pow"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0011" =>
                eclat_print_string(of_string("/"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0010" =>
                eclat_print_string(of_string("*"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0001" =>
                eclat_print_string(of_string("-"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when "0000" =>
                eclat_print_string(of_string("+"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              when others =>
                
              end case;
            when "0010" =>
              eclat_print_string(of_string("nil"));
              
              eclat_print_newline(eclat_unit);
              
              \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
              \state\ <= \$128_copy_args_to_heap544\;
            when "0001" =>
              \$764_n\ := \$v1651\(0 to 31);
              eclat_print_int(\$764_n\);
              
              eclat_print_newline(eclat_unit);
              
              \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
              \state\ <= \$128_copy_args_to_heap544\;
            when "0000" =>
              \$765_b\ := \$v1651\(0 to 0);
              \$v1655\ := \$765_b\;
              if \$v1655\(0) = '1' then
                eclat_print_string(of_string("true"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              else
                eclat_print_string(of_string("false"));
                
                eclat_print_newline(eclat_unit);
                
                \$128_copy_args_to_heap544_arg\ := eclat_sub(\$128_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$128_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$128_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                \state\ <= \$128_copy_args_to_heap544\;
              end if;
            when others =>
              
            end case;
          when pause_getII1667 =>
            \$arr1644_ptr_take\(0) := '0';
            \$769\ := \$arr1644_value\;
            \$v1665\ := \$arr1643_ptr_take\;
            if \$v1665\(0) = '1' then
              \state\ <= q_wait1664;
            else
              \$arr1643_ptr_take\(0) := '1';
              \$arr1643_ptr_write\ <= to_integer(unsigned(\$128_copy_args_to_heap544_arg\(64 to 95)));
              \$arr1643_write_request\ <= '1';
              \$arr1643_write\ <= \$769\;
              \state\ <= pause_setI1662;
            end if;
          when pause_getII1677 =>
            \$arr1644_ptr_take\(0) := '0';
            \$722\ := \$arr1644_value\;
            \$v1674\ := \$722\;
            \$v1675\ := \$v1674\(0 to 3);
            \$v1673\ := \$v1674\(4 to 67);
            case \$v1675\ is
            when "0001" =>
              \$723_a\ := \$v1673\(0 to 31);
              \$709_divisor\ := \$723_a\;
              \$v1672\ := eclat_eq(\$709_divisor\ & "00000000000000000000000000000000");
              if \$v1672\(0) = '1' then
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("Division par zero"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$718_forever5751608\;
              else
                \$130_div570_arg\ := eclat_sub(\$130_div570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$130_div570_arg\(32 to 63) & \$709_divisor\) & \$130_div570_arg\(64 to 95);
                \state\ <= \$130_div570\;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$727_forever5751609\;
            end case;
          when pause_getII1685 =>
            \$arr1644_ptr_take\(0) := '0';
            \$684_v\ := \$arr1644_value\;
            \$v1682\ := \$684_v\;
            \$v1683\ := \$v1682\(0 to 3);
            \$v1681\ := \$v1682\(4 to 67);
            case \$v1683\ is
            when "0001" =>
              \$690_a\ := \$v1681\(0 to 31);
              \$685_int_value\ := \$690_a\;
              \$131_mul571_arg\ := eclat_sub(\$131_mul571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$131_mul571_arg\(32 to 63) & \$685_int_value\) & \$131_mul571_arg\(64 to 95);
              \state\ <= \$131_mul571\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$694_forever5751610\;
            end case;
          when pause_getII1693 =>
            \$arr1644_ptr_take\(0) := '0';
            \$659_v\ := \$arr1644_value\;
            \$v1690\ := \$659_v\;
            \$v1691\ := \$v1690\(0 to 3);
            \$v1689\ := \$v1690\(4 to 67);
            case \$v1691\ is
            when "0001" =>
              \$665_a\ := \$v1689\(0 to 31);
              \$660_int_value\ := \$665_a\;
              \$132_sub572_arg\ := eclat_sub(\$132_sub572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$132_sub572_arg\(32 to 63) & \$660_int_value\) & \$132_sub572_arg\(64 to 95);
              \state\ <= \$132_sub572\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$669_forever5751611\;
            end case;
          when pause_getII1701 =>
            \$arr1644_ptr_take\(0) := '0';
            \$634_v\ := \$arr1644_value\;
            \$v1698\ := \$634_v\;
            \$v1699\ := \$v1698\(0 to 3);
            \$v1697\ := \$v1698\(4 to 67);
            case \$v1699\ is
            when "0001" =>
              \$640_a\ := \$v1697\(0 to 31);
              \$635_int_value\ := \$640_a\;
              \$133_add573_arg\ := eclat_sub(\$133_add573_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$133_add573_arg\(32 to 63) & \$635_int_value\) & \$133_add573_arg\(64 to 95);
              \state\ <= \$133_add573\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$644_forever5751612\;
            end case;
          when pause_setI1662 =>
            \$arr1643_write_request\ <= '0';
            \state\ <= pause_setII1663;
          when pause_setII1663 =>
            \$arr1643_ptr_take\(0) := '0';
            eclat_print_string(of_string("copy heap["));
            
            eclat_print_int(\$128_copy_args_to_heap544_arg\(64 to 95));
            
            eclat_print_string(of_string("] <-"));
            
            \$v1661\ := \$arr1644_ptr_take\;
            if \$v1661\(0) = '1' then
              \state\ <= q_wait1660;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$128_copy_args_to_heap544_arg\(32 to 63) & \$128_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI1658;
            end if;
          when q_wait1660 =>
            \$v1661\ := \$arr1644_ptr_take\;
            if \$v1661\(0) = '1' then
              \state\ <= q_wait1660;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$128_copy_args_to_heap544_arg\(32 to 63) & \$128_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI1658;
            end if;
          when q_wait1664 =>
            \$v1665\ := \$arr1643_ptr_take\;
            if \$v1665\(0) = '1' then
              \state\ <= q_wait1664;
            else
              \$arr1643_ptr_take\(0) := '1';
              \$arr1643_ptr_write\ <= to_integer(unsigned(\$128_copy_args_to_heap544_arg\(64 to 95)));
              \$arr1643_write_request\ <= '1';
              \$arr1643_write\ <= \$769\;
              \state\ <= pause_setI1662;
            end if;
          when q_wait1668 =>
            \$v1669\ := \$arr1644_ptr_take\;
            if \$v1669\(0) = '1' then
              \state\ <= q_wait1668;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$128_copy_args_to_heap544_arg\(32 to 63) & \$128_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI1666;
            end if;
          when q_wait1678 =>
            \$v1679\ := \$arr1644_ptr_take\;
            if \$v1679\(0) = '1' then
              \state\ <= q_wait1678;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_div570_arg\(0 to 31))));
              \state\ <= pause_getI1676;
            end if;
          when q_wait1686 =>
            \$v1687\ := \$arr1644_ptr_take\;
            if \$v1687\(0) = '1' then
              \state\ <= q_wait1686;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_mul571_arg\(0 to 31))));
              \state\ <= pause_getI1684;
            end if;
          when q_wait1694 =>
            \$v1695\ := \$arr1644_ptr_take\;
            if \$v1695\(0) = '1' then
              \state\ <= q_wait1694;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_sub572_arg\(0 to 31))));
              \state\ <= pause_getI1692;
            end if;
          when q_wait1702 =>
            \$v1703\ := \$arr1644_ptr_take\;
            if \$v1703\(0) = '1' then
              \state\ <= q_wait1702;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$133_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$133_add573_arg\(0 to 31))));
              \state\ <= pause_getI1700;
            end if;
          when compute1650 =>
            rdy1649 := eclat_false;
            case state_var2260 is
            when compute2110 =>
              rdy2109 := eclat_false;
              \$v2255\ := \$410\;
              if \$v2255\(0) = '1' then
                result2108 := eclat_true;
                rdy2109 := eclat_true;
                state_var2260 <= compute2110;
              else
                case state_var2261 is
                when \$415_copy_args_to_heap544\ =>
                  \$v2133\ := eclat_eq(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2133\(0) = '1' then
                    state_var2261 <= \$415_copy_args_to_heap544\;
                  else
                    \$v2132\ := \$arr1644_ptr_take\;
                    if \$v2132\(0) = '1' then
                      state_var2261 <= q_wait2131;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$415_copy_args_to_heap544_arg\(32 to 63) & \$415_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                      state_var2261 <= pause_getI2129;
                    end if;
                  end if;
                when \$416_pow569\ =>
                  \$v2134\ := eclat_eq(\$416_pow569_arg\(32 to 63) & "00000000000000000000000000000000");
                  if \$v2134\(0) = '1' then
                    state_var2261 <= \$416_pow569\;
                  else
                    \$416_pow569_arg\ := \$416_pow569_arg\(0 to 31) & eclat_sub(\$416_pow569_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$416_pow569_arg\(64 to 95) & \$416_pow569_arg\(0 to 31));
                    state_var2261 <= \$416_pow569\;
                  end if;
                when \$417_div570\ =>
                  \$v2143\ := eclat_eq(\$417_div570_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2143\(0) = '1' then
                    state_var2261 <= \$417_div570\;
                  else
                    \$v2142\ := \$arr1644_ptr_take\;
                    if \$v2142\(0) = '1' then
                      state_var2261 <= q_wait2141;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$417_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$417_div570_arg\(0 to 31))));
                      state_var2261 <= pause_getI2139;
                    end if;
                  end if;
                when \$418_mul571\ =>
                  \$v2151\ := eclat_eq(\$418_mul571_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2151\(0) = '1' then
                    state_var2261 <= \$418_mul571\;
                  else
                    \$v2150\ := \$arr1644_ptr_take\;
                    if \$v2150\(0) = '1' then
                      state_var2261 <= q_wait2149;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$418_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$418_mul571_arg\(0 to 31))));
                      state_var2261 <= pause_getI2147;
                    end if;
                  end if;
                when \$419_sub572\ =>
                  \$v2159\ := eclat_eq(\$419_sub572_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2159\(0) = '1' then
                    state_var2261 <= \$419_sub572\;
                  else
                    \$v2158\ := \$arr1644_ptr_take\;
                    if \$v2158\(0) = '1' then
                      state_var2261 <= q_wait2157;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$419_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$419_sub572_arg\(0 to 31))));
                      state_var2261 <= pause_getI2155;
                    end if;
                  end if;
                when \$420_add573\ =>
                  \$v2167\ := eclat_eq(\$420_add573_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2167\(0) = '1' then
                    state_var2261 <= \$420_add573\;
                  else
                    \$v2166\ := \$arr1644_ptr_take\;
                    if \$v2166\(0) = '1' then
                      state_var2261 <= q_wait2165;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$420_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$420_add573_arg\(0 to 31))));
                      state_var2261 <= pause_getI2163;
                    end if;
                  end if;
                when \$477_forever5751642\ =>
                  state_var2261 <= \$481_forever5751636\;
                when \$481_forever5751636\ =>
                  state_var2261 <= \$481_forever5751636\;
                when \$506_forever5751641\ =>
                  state_var2261 <= \$510_forever5751636\;
                when \$510_forever5751636\ =>
                  state_var2261 <= \$510_forever5751636\;
                when \$535_forever5751640\ =>
                  state_var2261 <= \$539_forever5751636\;
                when \$539_forever5751636\ =>
                  state_var2261 <= \$539_forever5751636\;
                when \$563_forever5751638\ =>
                  state_var2261 <= \$567_forever5751636\;
                when \$567_forever5751636\ =>
                  state_var2261 <= \$567_forever5751636\;
                when \$576_forever5751639\ =>
                  state_var2261 <= \$580_forever5751636\;
                when \$580_forever5751636\ =>
                  state_var2261 <= \$580_forever5751636\;
                when pause_getI2121 =>
                  state_var2261 <= pause_getII2122;
                when pause_getI2129 =>
                  state_var2261 <= pause_getII2130;
                when pause_getI2139 =>
                  state_var2261 <= pause_getII2140;
                when pause_getI2147 =>
                  state_var2261 <= pause_getII2148;
                when pause_getI2155 =>
                  state_var2261 <= pause_getII2156;
                when pause_getI2163 =>
                  state_var2261 <= pause_getII2164;
                when pause_getII2122 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$613\ := \$arr1644_value\;
                  \$v2119\ := \$613\;
                  \$v2120\ := \$v2119\(0 to 3);
                  \$v2114\ := \$v2119\(4 to 67);
                  case \$v2120\ is
                  when "0100" =>
                    eclat_print_string(of_string("fermeture"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                    state_var2261 <= \$415_copy_args_to_heap544\;
                  when "0011" =>
                    \$615_p\ := \$v2114\(0 to 4);
                    \$v2116\ := \$615_p\;
                    \$v2117\ := \$v2116\(0 to 3);
                    \$v2115\ := ""&\$v2116\(4);
                    case \$v2117\ is
                    when "0110" =>
                      eclat_print_string(of_string("<"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0101" =>
                      eclat_print_string(of_string("=="));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0100" =>
                      eclat_print_string(of_string("pow"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0011" =>
                      eclat_print_string(of_string("/"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0010" =>
                      eclat_print_string(of_string("*"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0001" =>
                      eclat_print_string(of_string("-"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when "0000" =>
                      eclat_print_string(of_string("+"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    when others =>
                      
                    end case;
                  when "0010" =>
                    eclat_print_string(of_string("nil"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                    state_var2261 <= \$415_copy_args_to_heap544\;
                  when "0001" =>
                    \$617_n\ := \$v2114\(0 to 31);
                    eclat_print_int(\$617_n\);
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                    state_var2261 <= \$415_copy_args_to_heap544\;
                  when "0000" =>
                    \$618_b\ := \$v2114\(0 to 0);
                    \$v2118\ := \$618_b\;
                    if \$v2118\(0) = '1' then
                      eclat_print_string(of_string("true"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    else
                      eclat_print_string(of_string("false"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$415_copy_args_to_heap544_arg\ := eclat_sub(\$415_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$415_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$415_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                      state_var2261 <= \$415_copy_args_to_heap544\;
                    end if;
                  when others =>
                    
                  end case;
                when pause_getII2130 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$622\ := \$arr1644_value\;
                  \$v2128\ := \$arr1643_ptr_take\;
                  if \$v2128\(0) = '1' then
                    state_var2261 <= q_wait2127;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr_write\ <= to_integer(unsigned(\$415_copy_args_to_heap544_arg\(64 to 95)));
                    \$arr1643_write_request\ <= '1';
                    \$arr1643_write\ <= \$622\;
                    state_var2261 <= pause_setI2125;
                  end if;
                when pause_getII2140 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$571\ := \$arr1644_value\;
                  \$v2137\ := \$571\;
                  \$v2138\ := \$v2137\(0 to 3);
                  \$v2136\ := \$v2137\(4 to 67);
                  case \$v2138\ is
                  when "0001" =>
                    \$572_a\ := \$v2136\(0 to 31);
                    \$554_divisor\ := \$572_a\;
                    \$v2135\ := eclat_eq(\$554_divisor\ & "00000000000000000000000000000000");
                    if \$v2135\(0) = '1' then
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("Division par zero"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var2261 <= \$563_forever5751638\;
                    else
                      \$417_div570_arg\ := eclat_sub(\$417_div570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$417_div570_arg\(32 to 63) & \$554_divisor\) & \$417_div570_arg\(64 to 95);
                      state_var2261 <= \$417_div570\;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2261 <= \$576_forever5751639\;
                  end case;
                when pause_getII2148 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$525_v\ := \$arr1644_value\;
                  \$v2145\ := \$525_v\;
                  \$v2146\ := \$v2145\(0 to 3);
                  \$v2144\ := \$v2145\(4 to 67);
                  case \$v2146\ is
                  when "0001" =>
                    \$531_a\ := \$v2144\(0 to 31);
                    \$526_int_value\ := \$531_a\;
                    \$418_mul571_arg\ := eclat_sub(\$418_mul571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$418_mul571_arg\(32 to 63) & \$526_int_value\) & \$418_mul571_arg\(64 to 95);
                    state_var2261 <= \$418_mul571\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2261 <= \$535_forever5751640\;
                  end case;
                when pause_getII2156 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$496_v\ := \$arr1644_value\;
                  \$v2153\ := \$496_v\;
                  \$v2154\ := \$v2153\(0 to 3);
                  \$v2152\ := \$v2153\(4 to 67);
                  case \$v2154\ is
                  when "0001" =>
                    \$502_a\ := \$v2152\(0 to 31);
                    \$497_int_value\ := \$502_a\;
                    \$419_sub572_arg\ := eclat_sub(\$419_sub572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$419_sub572_arg\(32 to 63) & \$497_int_value\) & \$419_sub572_arg\(64 to 95);
                    state_var2261 <= \$419_sub572\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2261 <= \$506_forever5751641\;
                  end case;
                when pause_getII2164 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$467_v\ := \$arr1644_value\;
                  \$v2161\ := \$467_v\;
                  \$v2162\ := \$v2161\(0 to 3);
                  \$v2160\ := \$v2161\(4 to 67);
                  case \$v2162\ is
                  when "0001" =>
                    \$473_a\ := \$v2160\(0 to 31);
                    \$468_int_value\ := \$473_a\;
                    \$420_add573_arg\ := eclat_sub(\$420_add573_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$420_add573_arg\(32 to 63) & \$468_int_value\) & \$420_add573_arg\(64 to 95);
                    state_var2261 <= \$420_add573\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2261 <= \$477_forever5751642\;
                  end case;
                when pause_setI2125 =>
                  \$arr1643_write_request\ <= '0';
                  state_var2261 <= pause_setII2126;
                when pause_setI2169 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2170;
                when pause_setI2174 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2175;
                when pause_setI2179 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2180;
                when pause_setI2185 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2186;
                when pause_setI2191 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2192;
                when pause_setI2196 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2197;
                when pause_setI2201 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2202;
                when pause_setI2206 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2207;
                when pause_setI2212 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2213;
                when pause_setI2217 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2218;
                when pause_setI2222 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2223;
                when pause_setI2229 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2230;
                when pause_setI2234 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2235;
                when pause_setI2239 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2240;
                when pause_setI2244 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2245;
                when pause_setI2249 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2261 <= pause_setII2250;
                when pause_setII2126 =>
                  \$arr1643_ptr_take\(0) := '0';
                  eclat_print_string(of_string("copy heap["));
                  
                  eclat_print_int(\$415_copy_args_to_heap544_arg\(64 to 95));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v2124\ := \$arr1644_ptr_take\;
                  if \$v2124\(0) = '1' then
                    state_var2261 <= q_wait2123;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$415_copy_args_to_heap544_arg\(32 to 63) & \$415_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var2261 <= pause_getI2121;
                  end if;
                when pause_setII2170 =>
                  \$arr1646_ptr_take\(0) := '0';
                  result2111 := eclat_unit;
                  rdy2112 := eclat_true;
                  state_var2261 <= compute2113;
                when pause_setII2175 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2172\ := \$arr1646_ptr_take\;
                  if \$v2172\(0) = '1' then
                    state_var2261 <= q_wait2171;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2168\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 15;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0111" & \$v2168\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2169;
                  end if;
                when pause_setII2180 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2177\ := \$arr1646_ptr_take\;
                  if \$v2177\(0) = '1' then
                    state_var2261 <= q_wait2176;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2173\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 14;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2173\&X"000000000";
                    state_var2261 <= pause_setI2174;
                  end if;
                when pause_setII2186 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2182\ := \$arr1646_ptr_take\;
                  if \$v2182\(0) = '1' then
                    state_var2261 <= q_wait2181;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2178\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 13;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0010" & \$v2178\&X"000000000";
                    state_var2261 <= pause_setI2179;
                  end if;
                when pause_setII2192 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2188\ := \$arr1646_ptr_take\;
                  if \$v2188\(0) = '1' then
                    state_var2261 <= q_wait2187;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2183\ := "00000000000000000000000000000001";
                    \$v2184\ := "0001" & \$v2183\&X"00000000";
                    \$arr1646_ptr_write\ <= 12;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2184\;
                    state_var2261 <= pause_setI2185;
                  end if;
                when pause_setII2197 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2194\ := \$arr1646_ptr_take\;
                  if \$v2194\(0) = '1' then
                    state_var2261 <= q_wait2193;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2189\ := "00000000000000000000000000000010";
                    \$v2190\ := "0001" & \$v2189\&X"00000000";
                    \$arr1646_ptr_write\ <= 11;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2190\;
                    state_var2261 <= pause_setI2191;
                  end if;
                when pause_setII2202 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2199\ := \$arr1646_ptr_take\;
                  if \$v2199\(0) = '1' then
                    state_var2261 <= q_wait2198;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2195\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 10;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0001" & \$v2195\&X"000000000";
                    state_var2261 <= pause_setI2196;
                  end if;
                when pause_setII2207 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2204\ := \$arr1646_ptr_take\;
                  if \$v2204\(0) = '1' then
                    state_var2261 <= q_wait2203;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2200\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 9;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0110" & \$v2200\&X"000000000";
                    state_var2261 <= pause_setI2201;
                  end if;
                when pause_setII2213 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2209\ := \$arr1646_ptr_take\;
                  if \$v2209\(0) = '1' then
                    state_var2261 <= q_wait2208;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2205\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 8;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2205\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2206;
                  end if;
                when pause_setII2218 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2215\ := \$arr1646_ptr_take\;
                  if \$v2215\(0) = '1' then
                    state_var2261 <= q_wait2214;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2210\ := eclat_unit;
                    \$v2211\ := "0010" & \$v2210\&"000"& X"000000000000000";
                    \$arr1646_ptr_write\ <= 7;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2211\;
                    state_var2261 <= pause_setI2212;
                  end if;
                when pause_setII2223 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2220\ := \$arr1646_ptr_take\;
                  if \$v2220\(0) = '1' then
                    state_var2261 <= q_wait2219;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2216\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 6;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2216\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2217;
                  end if;
                when pause_setII2230 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2225\ := \$arr1646_ptr_take\;
                  if \$v2225\(0) = '1' then
                    state_var2261 <= q_wait2224;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2221\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 5;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2221\&X"000000000";
                    state_var2261 <= pause_setI2222;
                  end if;
                when pause_setII2235 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2232\ := \$arr1646_ptr_take\;
                  if \$v2232\(0) = '1' then
                    state_var2261 <= q_wait2231;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2226\ := eclat_unit;
                    \$v2227\ := "0000" & \$v2226\;
                    \$v2228\ := "0011" & \$v2227\&"000"& X"00000000000000";
                    \$arr1646_ptr_write\ <= 4;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2228\;
                    state_var2261 <= pause_setI2229;
                  end if;
                when pause_setII2240 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2237\ := \$arr1646_ptr_take\;
                  if \$v2237\(0) = '1' then
                    state_var2261 <= q_wait2236;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2233\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 3;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2233\&X"000000000";
                    state_var2261 <= pause_setI2234;
                  end if;
                when pause_setII2245 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2242\ := \$arr1646_ptr_take\;
                  if \$v2242\(0) = '1' then
                    state_var2261 <= q_wait2241;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2238\ := "00000000000000000000000000000001";
                    \$arr1646_ptr_write\ <= 2;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2238\&X"000000000";
                    state_var2261 <= pause_setI2239;
                  end if;
                when pause_setII2250 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2247\ := \$arr1646_ptr_take\;
                  if \$v2247\(0) = '1' then
                    state_var2261 <= q_wait2246;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2243\ := "00000000000000000000000000001001";
                    \$arr1646_ptr_write\ <= 1;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1010" & \$v2243\&X"000000000";
                    state_var2261 <= pause_setI2244;
                  end if;
                when q_wait2123 =>
                  \$v2124\ := \$arr1644_ptr_take\;
                  if \$v2124\(0) = '1' then
                    state_var2261 <= q_wait2123;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$415_copy_args_to_heap544_arg\(32 to 63) & \$415_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var2261 <= pause_getI2121;
                  end if;
                when q_wait2127 =>
                  \$v2128\ := \$arr1643_ptr_take\;
                  if \$v2128\(0) = '1' then
                    state_var2261 <= q_wait2127;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr_write\ <= to_integer(unsigned(\$415_copy_args_to_heap544_arg\(64 to 95)));
                    \$arr1643_write_request\ <= '1';
                    \$arr1643_write\ <= \$622\;
                    state_var2261 <= pause_setI2125;
                  end if;
                when q_wait2131 =>
                  \$v2132\ := \$arr1644_ptr_take\;
                  if \$v2132\(0) = '1' then
                    state_var2261 <= q_wait2131;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$415_copy_args_to_heap544_arg\(32 to 63) & \$415_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var2261 <= pause_getI2129;
                  end if;
                when q_wait2141 =>
                  \$v2142\ := \$arr1644_ptr_take\;
                  if \$v2142\(0) = '1' then
                    state_var2261 <= q_wait2141;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$417_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$417_div570_arg\(0 to 31))));
                    state_var2261 <= pause_getI2139;
                  end if;
                when q_wait2149 =>
                  \$v2150\ := \$arr1644_ptr_take\;
                  if \$v2150\(0) = '1' then
                    state_var2261 <= q_wait2149;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$418_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$418_mul571_arg\(0 to 31))));
                    state_var2261 <= pause_getI2147;
                  end if;
                when q_wait2157 =>
                  \$v2158\ := \$arr1644_ptr_take\;
                  if \$v2158\(0) = '1' then
                    state_var2261 <= q_wait2157;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$419_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$419_sub572_arg\(0 to 31))));
                    state_var2261 <= pause_getI2155;
                  end if;
                when q_wait2165 =>
                  \$v2166\ := \$arr1644_ptr_take\;
                  if \$v2166\(0) = '1' then
                    state_var2261 <= q_wait2165;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$420_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$420_add573_arg\(0 to 31))));
                    state_var2261 <= pause_getI2163;
                  end if;
                when q_wait2171 =>
                  \$v2172\ := \$arr1646_ptr_take\;
                  if \$v2172\(0) = '1' then
                    state_var2261 <= q_wait2171;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2168\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 15;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0111" & \$v2168\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2169;
                  end if;
                when q_wait2176 =>
                  \$v2177\ := \$arr1646_ptr_take\;
                  if \$v2177\(0) = '1' then
                    state_var2261 <= q_wait2176;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2173\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 14;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2173\&X"000000000";
                    state_var2261 <= pause_setI2174;
                  end if;
                when q_wait2181 =>
                  \$v2182\ := \$arr1646_ptr_take\;
                  if \$v2182\(0) = '1' then
                    state_var2261 <= q_wait2181;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2178\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 13;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0010" & \$v2178\&X"000000000";
                    state_var2261 <= pause_setI2179;
                  end if;
                when q_wait2187 =>
                  \$v2188\ := \$arr1646_ptr_take\;
                  if \$v2188\(0) = '1' then
                    state_var2261 <= q_wait2187;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2183\ := "00000000000000000000000000000001";
                    \$v2184\ := "0001" & \$v2183\&X"00000000";
                    \$arr1646_ptr_write\ <= 12;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2184\;
                    state_var2261 <= pause_setI2185;
                  end if;
                when q_wait2193 =>
                  \$v2194\ := \$arr1646_ptr_take\;
                  if \$v2194\(0) = '1' then
                    state_var2261 <= q_wait2193;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2189\ := "00000000000000000000000000000010";
                    \$v2190\ := "0001" & \$v2189\&X"00000000";
                    \$arr1646_ptr_write\ <= 11;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2190\;
                    state_var2261 <= pause_setI2191;
                  end if;
                when q_wait2198 =>
                  \$v2199\ := \$arr1646_ptr_take\;
                  if \$v2199\(0) = '1' then
                    state_var2261 <= q_wait2198;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2195\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 10;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0001" & \$v2195\&X"000000000";
                    state_var2261 <= pause_setI2196;
                  end if;
                when q_wait2203 =>
                  \$v2204\ := \$arr1646_ptr_take\;
                  if \$v2204\(0) = '1' then
                    state_var2261 <= q_wait2203;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2200\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 9;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0110" & \$v2200\&X"000000000";
                    state_var2261 <= pause_setI2201;
                  end if;
                when q_wait2208 =>
                  \$v2209\ := \$arr1646_ptr_take\;
                  if \$v2209\(0) = '1' then
                    state_var2261 <= q_wait2208;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2205\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 8;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2205\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2206;
                  end if;
                when q_wait2214 =>
                  \$v2215\ := \$arr1646_ptr_take\;
                  if \$v2215\(0) = '1' then
                    state_var2261 <= q_wait2214;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2210\ := eclat_unit;
                    \$v2211\ := "0010" & \$v2210\&"000"& X"000000000000000";
                    \$arr1646_ptr_write\ <= 7;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2211\;
                    state_var2261 <= pause_setI2212;
                  end if;
                when q_wait2219 =>
                  \$v2220\ := \$arr1646_ptr_take\;
                  if \$v2220\(0) = '1' then
                    state_var2261 <= q_wait2219;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2216\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 6;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2216\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2217;
                  end if;
                when q_wait2224 =>
                  \$v2225\ := \$arr1646_ptr_take\;
                  if \$v2225\(0) = '1' then
                    state_var2261 <= q_wait2224;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2221\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 5;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2221\&X"000000000";
                    state_var2261 <= pause_setI2222;
                  end if;
                when q_wait2231 =>
                  \$v2232\ := \$arr1646_ptr_take\;
                  if \$v2232\(0) = '1' then
                    state_var2261 <= q_wait2231;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2226\ := eclat_unit;
                    \$v2227\ := "0000" & \$v2226\;
                    \$v2228\ := "0011" & \$v2227\&"000"& X"00000000000000";
                    \$arr1646_ptr_write\ <= 4;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2228\;
                    state_var2261 <= pause_setI2229;
                  end if;
                when q_wait2236 =>
                  \$v2237\ := \$arr1646_ptr_take\;
                  if \$v2237\(0) = '1' then
                    state_var2261 <= q_wait2236;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2233\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 3;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2233\&X"000000000";
                    state_var2261 <= pause_setI2234;
                  end if;
                when q_wait2241 =>
                  \$v2242\ := \$arr1646_ptr_take\;
                  if \$v2242\(0) = '1' then
                    state_var2261 <= q_wait2241;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2238\ := "00000000000000000000000000000001";
                    \$arr1646_ptr_write\ <= 2;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2238\&X"000000000";
                    state_var2261 <= pause_setI2239;
                  end if;
                when q_wait2246 =>
                  \$v2247\ := \$arr1646_ptr_take\;
                  if \$v2247\(0) = '1' then
                    state_var2261 <= q_wait2246;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2243\ := "00000000000000000000000000001001";
                    \$arr1646_ptr_write\ <= 1;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1010" & \$v2243\&X"000000000";
                    state_var2261 <= pause_setI2244;
                  end if;
                when q_wait2251 =>
                  \$v2252\ := \$arr1646_ptr_take\;
                  if \$v2252\(0) = '1' then
                    state_var2261 <= q_wait2251;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2248\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 0;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0000" & \$v2248\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2249;
                  end if;
                when compute2113 =>
                  rdy2112 := eclat_false;
                  \$v2252\ := \$arr1646_ptr_take\;
                  if \$v2252\(0) = '1' then
                    state_var2261 <= q_wait2251;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2248\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 0;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0000" & \$v2248\&"000"& X"0000000000000000";
                    state_var2261 <= pause_setI2249;
                  end if;
                end case;
                \$v2254\ := eclat_not(rdy2112);
                if \$v2254\(0) = '1' then
                  result2111 := eclat_unit;
                end if;
                \$412\ := result2111 & rdy2112;
                result2108 := ""&\$412\(1);
                rdy2109 := eclat_true;
                state_var2260 <= compute2110;
              end if;
            end case;
            \$v2257\ := eclat_not(rdy2109);
            if \$v2257\(0) = '1' then
              result2108 := eclat_false;
            end if;
            \$410\ := result2108;
            \$135_is_loaded\ := result2108;
            case state_var2259 is
            when compute2105 =>
              rdy2104 := eclat_false;
              result2103 := eclat_if(\$135_is_loaded\ & eclat_add(\$408\ & "00000000000000000000000000000001") & \$408\);
              rdy2104 := eclat_true;
              state_var2259 <= compute2105;
            end case;
            \$v2107\ := eclat_not(rdy2104);
            if \$v2107\(0) = '1' then
              result2103 := "00000000000000000000000000000000";
            end if;
            \$408\ := result2103;
            \$136_cy\ := result2103;
            case state_var2258 is
            when \$118_forever5741614\ =>
              state_var2258 <= \$118_forever5741614\;
            when \$118_forever5741621\ =>
              state_var2258 <= \$118_forever5741614\;
            when \$118_forever5741622\ =>
              state_var2258 <= \$118_forever5741614\;
            when \$118_forever5741623\ =>
              state_var2258 <= \$118_forever5741614\;
            when \$118_forever5741624\ =>
              state_var2258 <= \$118_forever5741614\;
            when \$121_forever5751613\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751625\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751626\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751627\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751628\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751629\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751630\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751631\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751632\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751633\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751634\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$121_forever5751635\ =>
              state_var2258 <= \$121_forever5751613\;
            when \$144_copy_args_to_heap544\ =>
              \$v1728\ := eclat_eq(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1728\(0) = '1' then
                \$144_copy_args_to_heap544_result\ := \$144_copy_args_to_heap544_arg\(32 to 63);
                \$v1773\ := \$arr1647_ptr_take\;
                if \$v1773\(0) = '1' then
                  state_var2258 <= q_wait1772;
                else
                  \$arr1647_ptr_take\(0) := '1';
                  \$arr1647_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(96 to 127)));
                  \$arr1647_write_request\ <= '1';
                  \$arr1647_write\ <= eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127);
                  state_var2258 <= pause_setI1770;
                end if;
              else
                \$v1727\ := \$arr1644_ptr_take\;
                if \$v1727\(0) = '1' then
                  state_var2258 <= q_wait1726;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$144_copy_args_to_heap544_arg\(32 to 63) & \$144_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1724;
                end if;
              end if;
            when \$145_pow569\ =>
              \$v1729\ := eclat_eq(\$145_pow569_arg\(32 to 63) & "00000000000000000000000000000000");
              if \$v1729\(0) = '1' then
                \$145_pow569_result\ := \$145_pow569_arg\(64 to 95);
                resultat := \$145_pow569_result\;
                \$v1869\ := \$arr1644_ptr_take\;
                if \$v1869\(0) = '1' then
                  state_var2258 <= q_wait1868;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1866;
                end if;
              else
                \$145_pow569_arg\ := \$145_pow569_arg\(0 to 31) & eclat_sub(\$145_pow569_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$145_pow569_arg\(64 to 95) & \$145_pow569_arg\(0 to 31));
                state_var2258 <= \$145_pow569\;
              end if;
            when \$146_div570\ =>
              \$v1738\ := eclat_eq(\$146_div570_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1738\(0) = '1' then
                \$146_div570_result\ := \$146_div570_arg\(32 to 63);
                resultat := \$146_div570_result\;
                \$v1888\ := \$arr1644_ptr_take\;
                if \$v1888\(0) = '1' then
                  state_var2258 <= q_wait1887;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1885;
                end if;
              else
                \$v1737\ := \$arr1644_ptr_take\;
                if \$v1737\(0) = '1' then
                  state_var2258 <= q_wait1736;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_div570_arg\(0 to 31))));
                  state_var2258 <= pause_getI1734;
                end if;
              end if;
            when \$147_mul571\ =>
              \$v1746\ := eclat_eq(\$147_mul571_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1746\(0) = '1' then
                \$147_mul571_result\ := \$147_mul571_arg\(32 to 63);
                resultat := \$147_mul571_result\;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1933\ := \$arr1644_ptr_take\;
                if \$v1933\(0) = '1' then
                  state_var2258 <= q_wait1932;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1930;
                end if;
              else
                \$v1745\ := \$arr1644_ptr_take\;
                if \$v1745\(0) = '1' then
                  state_var2258 <= q_wait1744;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_mul571_arg\(0 to 31))));
                  state_var2258 <= pause_getI1742;
                end if;
              end if;
            when \$148_sub572\ =>
              \$v1754\ := eclat_eq(\$148_sub572_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1754\(0) = '1' then
                \$148_sub572_result\ := \$148_sub572_arg\(32 to 63);
                resultat := \$148_sub572_result\;
                \$v1949\ := \$arr1644_ptr_take\;
                if \$v1949\(0) = '1' then
                  state_var2258 <= q_wait1948;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1945\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & \$v1945\&X"00000000";
                  state_var2258 <= pause_setI1946;
                end if;
              else
                \$v1753\ := \$arr1644_ptr_take\;
                if \$v1753\(0) = '1' then
                  state_var2258 <= q_wait1752;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_sub572_arg\(0 to 31))));
                  state_var2258 <= pause_getI1750;
                end if;
              end if;
            when \$149_add573\ =>
              \$v1762\ := eclat_eq(\$149_add573_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1762\(0) = '1' then
                \$149_add573_result\ := \$149_add573_arg\(32 to 63);
                resultat := \$149_add573_result\;
                \$v1994\ := \$arr1644_ptr_take\;
                if \$v1994\(0) = '1' then
                  state_var2258 <= q_wait1993;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1991;
                end if;
              else
                \$v1761\ := \$arr1644_ptr_take\;
                if \$v1761\(0) = '1' then
                  state_var2258 <= q_wait1760;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$149_add573_arg\(0 to 31))));
                  state_var2258 <= pause_getI1758;
                end if;
              end if;
            when \$150_vm_run_code547\ =>
              \$v2099\ := ""&\$150_vm_run_code547_arg\(294);
              if \$v2099\(0) = '1' then
                eclat_print_string(of_string("[sp:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(0 to 31));
                
                eclat_print_string(of_string("|env:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(32 to 63));
                
                eclat_print_string(of_string("|pc:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(64 to 95));
                
                eclat_print_string(of_string("|fp:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(96 to 127));
                
                eclat_print_string(of_string("]"));
                
                eclat_print_string(of_string("|gp:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(128 to 159));
                
                eclat_print_string(of_string("|hp:"));
                
                eclat_print_int(\$150_vm_run_code547_arg\(128 to 159));
                
                eclat_print_newline(eclat_unit);
                
                \$v2098\ := \$arr1646_ptr_take\;
                if \$v2098\(0) = '1' then
                  state_var2258 <= q_wait2097;
                else
                  \$arr1646_ptr_take\(0) := '1';
                  \$arr1646_ptr\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(64 to 95)));
                  state_var2258 <= pause_getI2095;
                end if;
              else
                \$v2098\ := \$arr1646_ptr_take\;
                if \$v2098\(0) = '1' then
                  state_var2258 <= q_wait2097;
                else
                  \$arr1646_ptr_take\(0) := '1';
                  \$arr1646_ptr\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(64 to 95)));
                  state_var2258 <= pause_getI2095;
                end if;
              end if;
            when \$209_forever5741620\ =>
              state_var2258 <= \$213_forever5741614\;
            when \$213_forever5741614\ =>
              state_var2258 <= \$213_forever5741614\;
            when \$259_forever5751619\ =>
              state_var2258 <= \$263_forever5751613\;
            when \$263_forever5751613\ =>
              state_var2258 <= \$263_forever5751613\;
            when \$288_forever5751618\ =>
              state_var2258 <= \$292_forever5751613\;
            when \$292_forever5751613\ =>
              state_var2258 <= \$292_forever5751613\;
            when \$317_forever5751617\ =>
              state_var2258 <= \$321_forever5751613\;
            when \$321_forever5751613\ =>
              state_var2258 <= \$321_forever5751613\;
            when \$345_forever5751615\ =>
              state_var2258 <= \$349_forever5751613\;
            when \$349_forever5751613\ =>
              state_var2258 <= \$349_forever5751613\;
            when \$358_forever5751616\ =>
              state_var2258 <= \$362_forever5751613\;
            when \$362_forever5751613\ =>
              state_var2258 <= \$362_forever5751613\;
            when pause_getI1716 =>
              state_var2258 <= pause_getII1717;
            when pause_getI1724 =>
              state_var2258 <= pause_getII1725;
            when pause_getI1734 =>
              state_var2258 <= pause_getII1735;
            when pause_getI1742 =>
              state_var2258 <= pause_getII1743;
            when pause_getI1750 =>
              state_var2258 <= pause_getII1751;
            when pause_getI1758 =>
              state_var2258 <= pause_getII1759;
            when pause_getI1796 =>
              state_var2258 <= pause_getII1797;
            when pause_getI1800 =>
              state_var2258 <= pause_getII1801;
            when pause_getI1825 =>
              state_var2258 <= pause_getII1826;
            when pause_getI1836 =>
              state_var2258 <= pause_getII1837;
            when pause_getI1847 =>
              state_var2258 <= pause_getII1848;
            when pause_getI1854 =>
              state_var2258 <= pause_getII1855;
            when pause_getI1861 =>
              state_var2258 <= pause_getII1862;
            when pause_getI1873 =>
              state_var2258 <= pause_getII1874;
            when pause_getI1880 =>
              state_var2258 <= pause_getII1881;
            when pause_getI1892 =>
              state_var2258 <= pause_getII1893;
            when pause_getI1908 =>
              state_var2258 <= pause_getII1909;
            when pause_getI1919 =>
              state_var2258 <= pause_getII1920;
            when pause_getI1930 =>
              state_var2258 <= pause_getII1931;
            when pause_getI1941 =>
              state_var2258 <= pause_getII1942;
            when pause_getI1957 =>
              state_var2258 <= pause_getII1958;
            when pause_getI1968 =>
              state_var2258 <= pause_getII1969;
            when pause_getI1979 =>
              state_var2258 <= pause_getII1980;
            when pause_getI1986 =>
              state_var2258 <= pause_getII1987;
            when pause_getI1999 =>
              state_var2258 <= pause_getII2000;
            when pause_getI2012 =>
              state_var2258 <= pause_getII2013;
            when pause_getI2016 =>
              state_var2258 <= pause_getII2017;
            when pause_getI2023 =>
              state_var2258 <= pause_getII2024;
            when pause_getI2030 =>
              state_var2258 <= pause_getII2031;
            when pause_getI2038 =>
              state_var2258 <= pause_getII2039;
            when pause_getI2046 =>
              state_var2258 <= pause_getII2047;
            when pause_getI2057 =>
              state_var2258 <= pause_getII2058;
            when pause_getI2065 =>
              state_var2258 <= pause_getII2066;
            when pause_getI2073 =>
              state_var2258 <= pause_getII2074;
            when pause_getI2084 =>
              state_var2258 <= pause_getII2085;
            when pause_getI2095 =>
              state_var2258 <= pause_getII2096;
            when pause_getII1717 =>
              \$arr1644_ptr_take\(0) := '0';
              \$395\ := \$arr1644_value\;
              \$v1714\ := \$395\;
              \$v1715\ := \$v1714\(0 to 3);
              \$v1709\ := \$v1714\(4 to 67);
              case \$v1715\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                state_var2258 <= \$144_copy_args_to_heap544\;
              when "0011" =>
                \$397_p\ := \$v1709\(0 to 4);
                \$v1711\ := \$397_p\;
                \$v1712\ := \$v1711\(0 to 3);
                \$v1710\ := ""&\$v1711\(4);
                case \$v1712\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                state_var2258 <= \$144_copy_args_to_heap544\;
              when "0001" =>
                \$399_n\ := \$v1709\(0 to 31);
                eclat_print_int(\$399_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                state_var2258 <= \$144_copy_args_to_heap544\;
              when "0000" =>
                \$400_b\ := \$v1709\(0 to 0);
                \$v1713\ := \$400_b\;
                if \$v1713\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$144_copy_args_to_heap544_arg\ := eclat_sub(\$144_copy_args_to_heap544_arg\(0 to 31) & "00000000000000000000000000000001") & \$144_copy_args_to_heap544_arg\(32 to 63) & eclat_add(\$144_copy_args_to_heap544_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2258 <= \$144_copy_args_to_heap544\;
                end if;
              when others =>
                
              end case;
            when pause_getII1725 =>
              \$arr1644_ptr_take\(0) := '0';
              \$404\ := \$arr1644_value\;
              \$v1723\ := \$arr1643_ptr_take\;
              if \$v1723\(0) = '1' then
                state_var2258 <= q_wait1722;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(\$144_copy_args_to_heap544_arg\(64 to 95)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= \$404\;
                state_var2258 <= pause_setI1720;
              end if;
            when pause_getII1735 =>
              \$arr1644_ptr_take\(0) := '0';
              \$353\ := \$arr1644_value\;
              \$v1732\ := \$353\;
              \$v1733\ := \$v1732\(0 to 3);
              \$v1731\ := \$v1732\(4 to 67);
              case \$v1733\ is
              when "0001" =>
                \$354_a\ := \$v1731\(0 to 31);
                \$336_divisor\ := \$354_a\;
                \$v1730\ := eclat_eq(\$336_divisor\ & "00000000000000000000000000000000");
                if \$v1730\(0) = '1' then
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("Division par zero"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2258 <= \$345_forever5751615\;
                else
                  \$146_div570_arg\ := eclat_sub(\$146_div570_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$146_div570_arg\(32 to 63) & \$336_divisor\) & \$146_div570_arg\(64 to 95);
                  state_var2258 <= \$146_div570\;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$358_forever5751616\;
              end case;
            when pause_getII1743 =>
              \$arr1644_ptr_take\(0) := '0';
              \$307_v\ := \$arr1644_value\;
              \$v1740\ := \$307_v\;
              \$v1741\ := \$v1740\(0 to 3);
              \$v1739\ := \$v1740\(4 to 67);
              case \$v1741\ is
              when "0001" =>
                \$313_a\ := \$v1739\(0 to 31);
                \$308_int_value\ := \$313_a\;
                \$147_mul571_arg\ := eclat_sub(\$147_mul571_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$147_mul571_arg\(32 to 63) & \$308_int_value\) & \$147_mul571_arg\(64 to 95);
                state_var2258 <= \$147_mul571\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$317_forever5751617\;
              end case;
            when pause_getII1751 =>
              \$arr1644_ptr_take\(0) := '0';
              \$278_v\ := \$arr1644_value\;
              \$v1748\ := \$278_v\;
              \$v1749\ := \$v1748\(0 to 3);
              \$v1747\ := \$v1748\(4 to 67);
              case \$v1749\ is
              when "0001" =>
                \$284_a\ := \$v1747\(0 to 31);
                \$279_int_value\ := \$284_a\;
                \$148_sub572_arg\ := eclat_sub(\$148_sub572_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$148_sub572_arg\(32 to 63) & \$279_int_value\) & \$148_sub572_arg\(64 to 95);
                state_var2258 <= \$148_sub572\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$288_forever5751618\;
              end case;
            when pause_getII1759 =>
              \$arr1644_ptr_take\(0) := '0';
              \$249_v\ := \$arr1644_value\;
              \$v1756\ := \$249_v\;
              \$v1757\ := \$v1756\(0 to 3);
              \$v1755\ := \$v1756\(4 to 67);
              case \$v1757\ is
              when "0001" =>
                \$255_a\ := \$v1755\(0 to 31);
                \$250_int_value\ := \$255_a\;
                \$149_add573_arg\ := eclat_sub(\$149_add573_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$149_add573_arg\(32 to 63) & \$250_int_value\) & \$149_add573_arg\(64 to 95);
                state_var2258 <= \$149_add573\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$259_forever5751619\;
              end case;
            when pause_getII1797 =>
              \$arr1644_ptr_take\(0) := '0';
              second_value := \$arr1644_value\;
              \$v1794\ := first_value;
              \$v1795\ := \$v1794\(0 to 3);
              \$v1784\ := \$v1794\(4 to 67);
              case \$v1795\ is
              when "0010" =>
                \$v1786\ := second_value;
                \$v1787\ := \$v1786\(0 to 3);
                \$v1785\ := \$v1786\(4 to 67);
                case \$v1787\ is
                when "0010" =>
                  res := eclat_true;
                  \$v1783\ := \$arr1644_ptr_take\;
                  if \$v1783\(0) = '1' then
                    state_var2258 <= q_wait1782;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$193_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1780;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2258 <= \$118_forever5741622\;
                end case;
              when "0000" =>
                \$99_a1\ := \$v1784\(0 to 0);
                \$v1789\ := second_value;
                \$v1790\ := \$v1789\(0 to 3);
                \$v1788\ := \$v1789\(4 to 67);
                case \$v1790\ is
                when "0000" =>
                  b2 := \$v1788\(0 to 0);
                  res := eclat_if(\$99_a1\ & eclat_if(b2 & eclat_true & eclat_false) & 
                         eclat_if(b2 & eclat_false & eclat_true));
                  \$v1783\ := \$arr1644_ptr_take\;
                  if \$v1783\(0) = '1' then
                    state_var2258 <= q_wait1782;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$193_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1780;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2258 <= \$118_forever5741623\;
                end case;
              when "0001" =>
                \$100_a\ := \$v1784\(0 to 31);
                \$v1792\ := second_value;
                \$v1793\ := \$v1792\(0 to 3);
                \$v1791\ := \$v1792\(4 to 67);
                case \$v1793\ is
                when "0001" =>
                  b := \$v1791\(0 to 31);
                  res := eclat_eq(\$100_a\ & b);
                  \$v1783\ := \$arr1644_ptr_take\;
                  if \$v1783\(0) = '1' then
                    state_var2258 <= q_wait1782;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$193_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1780;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2258 <= \$118_forever5741624\;
                end case;
              when others =>
                eclat_print_string(of_string("il n'y a pas d'égalité possible \n"));
                
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$118_forever5741621\;
              end case;
            when pause_getII1801 =>
              \$arr1644_ptr_take\(0) := '0';
              first_value := \$arr1644_value\;
              \$v1799\ := \$arr1644_ptr_take\;
              if \$v1799\(0) = '1' then
                state_var2258 <= q_wait1798;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2258 <= pause_getI1796;
              end if;
            when pause_getII1826 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v57\ := \$arr1644_value\;
              \$v1823\ := \$v57\;
              \$v1824\ := \$v1823\(0 to 3);
              \$v1818\ := \$v1823\(4 to 67);
              case \$v1824\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2258 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1813\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                  state_var2258 <= pause_setI1814;
                end if;
              when "0011" =>
                \$114_p\ := \$v1818\(0 to 4);
                \$v1820\ := \$114_p\;
                \$v1821\ := \$v1820\(0 to 3);
                \$v1819\ := ""&\$v1820\(4);
                case \$v1821\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2258 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1813\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                  state_var2258 <= pause_setI1814;
                end if;
              when "0001" =>
                \$115_n\ := \$v1818\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2258 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1813\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                  state_var2258 <= pause_setI1814;
                end if;
              when "0000" =>
                \$116_b\ := \$v1818\(0 to 0);
                \$v1822\ := \$116_b\;
                if \$v1822\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2258 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1813\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                    state_var2258 <= pause_setI1814;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1837 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v54\ := \$arr1644_value\;
              \$v1834\ := \$v54\;
              \$v1835\ := \$v1834\(0 to 3);
              \$v1829\ := \$v1834\(4 to 67);
              case \$v1835\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1828\ := \$arr1644_ptr_take\;
                if \$v1828\(0) = '1' then
                  state_var2258 <= q_wait1827;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1825;
                end if;
              when "0011" =>
                \$114_p\ := \$v1829\(0 to 4);
                \$v1831\ := \$114_p\;
                \$v1832\ := \$v1831\(0 to 3);
                \$v1830\ := ""&\$v1831\(4);
                case \$v1832\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1828\ := \$arr1644_ptr_take\;
                if \$v1828\(0) = '1' then
                  state_var2258 <= q_wait1827;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1825;
                end if;
              when "0001" =>
                \$115_n\ := \$v1829\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1828\ := \$arr1644_ptr_take\;
                if \$v1828\(0) = '1' then
                  state_var2258 <= q_wait1827;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1825;
                end if;
              when "0000" =>
                \$116_b\ := \$v1829\(0 to 0);
                \$v1833\ := \$116_b\;
                if \$v1833\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1828\ := \$arr1644_ptr_take\;
                  if \$v1828\(0) = '1' then
                    state_var2258 <= q_wait1827;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1825;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1848 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v51\ := \$arr1644_value\;
              \$v1845\ := \$v51\;
              \$v1846\ := \$v1845\(0 to 3);
              \$v1840\ := \$v1845\(4 to 67);
              case \$v1846\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1839\ := \$arr1644_ptr_take\;
                if \$v1839\(0) = '1' then
                  state_var2258 <= q_wait1838;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2258 <= pause_getI1836;
                end if;
              when "0011" =>
                \$114_p\ := \$v1840\(0 to 4);
                \$v1842\ := \$114_p\;
                \$v1843\ := \$v1842\(0 to 3);
                \$v1841\ := ""&\$v1842\(4);
                case \$v1843\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1839\ := \$arr1644_ptr_take\;
                if \$v1839\(0) = '1' then
                  state_var2258 <= q_wait1838;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2258 <= pause_getI1836;
                end if;
              when "0001" =>
                \$115_n\ := \$v1840\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1839\ := \$arr1644_ptr_take\;
                if \$v1839\(0) = '1' then
                  state_var2258 <= q_wait1838;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2258 <= pause_getI1836;
                end if;
              when "0000" =>
                \$116_b\ := \$v1840\(0 to 0);
                \$v1844\ := \$116_b\;
                if \$v1844\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1839\ := \$arr1644_ptr_take\;
                  if \$v1839\(0) = '1' then
                    state_var2258 <= q_wait1838;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2258 <= pause_getI1836;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1855 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v48\ := \$arr1644_value\;
              \$v1852\ := \$v48\;
              \$v1853\ := \$v1852\(0 to 3);
              \$v1851\ := \$v1852\(4 to 67);
              case \$v1853\ is
              when "0001" =>
                a := \$v1851\(0 to 31);
                scd_operand := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1850\ := \$arr1644_ptr_take\;
                if \$v1850\(0) = '1' then
                  state_var2258 <= q_wait1849;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                  state_var2258 <= pause_getI1847;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751626\;
              end case;
            when pause_getII1862 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v46\ := \$arr1644_value\;
              \$v1859\ := \$v46\;
              \$v1860\ := \$v1859\(0 to 3);
              \$v1858\ := \$v1859\(4 to 67);
              case \$v1860\ is
              when "0001" =>
                a := \$v1858\(0 to 31);
                fst_operand := a;
                \$v1857\ := \$arr1644_ptr_take\;
                if \$v1857\(0) = '1' then
                  state_var2258 <= q_wait1856;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2258 <= pause_getI1854;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751627\;
              end case;
            when pause_getII1874 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v69\ := \$arr1644_value\;
              \$v1871\ := \$v69\;
              \$v1872\ := \$v1871\(0 to 3);
              \$v1870\ := \$v1871\(4 to 67);
              case \$v1872\ is
              when "0001" =>
                a := \$v1870\(0 to 31);
                exponent := a;
                \$145_pow569_arg\ := base & exponent & "00000000000000000000000000000001";
                state_var2258 <= \$145_pow569\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751629\;
              end case;
            when pause_getII1881 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v67\ := \$arr1644_value\;
              \$v1878\ := \$v67\;
              \$v1879\ := \$v1878\(0 to 3);
              \$v1877\ := \$v1878\(4 to 67);
              case \$v1879\ is
              when "0001" =>
                a := \$v1877\(0 to 31);
                base := a;
                \$v1876\ := \$arr1644_ptr_take\;
                if \$v1876\(0) = '1' then
                  state_var2258 <= q_wait1875;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2258 <= pause_getI1873;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751630\;
              end case;
            when pause_getII1893 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v93\ := \$arr1644_value\;
              \$v1890\ := \$v93\;
              \$v1891\ := \$v1890\(0 to 3);
              \$v1889\ := \$v1890\(4 to 67);
              case \$v1891\ is
              when "0001" =>
                a := \$v1889\(0 to 31);
                debut := a;
                \$146_div570_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                state_var2258 <= \$146_div570\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751632\;
              end case;
            when pause_getII1909 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v125\ := \$arr1644_value\;
              \$v1906\ := \$v125\;
              \$v1907\ := \$v1906\(0 to 3);
              \$v1901\ := \$v1906\(4 to 67);
              case \$v1907\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2258 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1897;
                end if;
              when "0011" =>
                \$114_p\ := \$v1901\(0 to 4);
                \$v1903\ := \$114_p\;
                \$v1904\ := \$v1903\(0 to 3);
                \$v1902\ := ""&\$v1903\(4);
                case \$v1904\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2258 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1897;
                end if;
              when "0001" =>
                \$115_n\ := \$v1901\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2258 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2258 <= pause_setI1897;
                end if;
              when "0000" =>
                \$116_b\ := \$v1901\(0 to 0);
                \$v1905\ := \$116_b\;
                if \$v1905\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2258 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2258 <= pause_setI1897;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1920 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v118\ := \$arr1644_value\;
              \$v1917\ := \$v118\;
              \$v1918\ := \$v1917\(0 to 3);
              \$v1912\ := \$v1917\(4 to 67);
              case \$v1918\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1911\ := \$arr1644_ptr_take\;
                if \$v1911\(0) = '1' then
                  state_var2258 <= q_wait1910;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1908;
                end if;
              when "0011" =>
                \$114_p\ := \$v1912\(0 to 4);
                \$v1914\ := \$114_p\;
                \$v1915\ := \$v1914\(0 to 3);
                \$v1913\ := ""&\$v1914\(4);
                case \$v1915\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1911\ := \$arr1644_ptr_take\;
                if \$v1911\(0) = '1' then
                  state_var2258 <= q_wait1910;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1908;
                end if;
              when "0001" =>
                \$115_n\ := \$v1912\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1911\ := \$arr1644_ptr_take\;
                if \$v1911\(0) = '1' then
                  state_var2258 <= q_wait1910;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1908;
                end if;
              when "0000" =>
                \$116_b\ := \$v1912\(0 to 0);
                \$v1916\ := \$116_b\;
                if \$v1916\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1911\ := \$arr1644_ptr_take\;
                  if \$v1911\(0) = '1' then
                    state_var2258 <= q_wait1910;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1908;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1931 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v115\ := \$arr1644_value\;
              \$v1928\ := \$v115\;
              \$v1929\ := \$v1928\(0 to 3);
              \$v1923\ := \$v1928\(4 to 67);
              case \$v1929\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1922\ := \$arr1644_ptr_take\;
                if \$v1922\(0) = '1' then
                  state_var2258 <= q_wait1921;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1919;
                end if;
              when "0011" =>
                \$114_p\ := \$v1923\(0 to 4);
                \$v1925\ := \$114_p\;
                \$v1926\ := \$v1925\(0 to 3);
                \$v1924\ := ""&\$v1925\(4);
                case \$v1926\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1922\ := \$arr1644_ptr_take\;
                if \$v1922\(0) = '1' then
                  state_var2258 <= q_wait1921;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1919;
                end if;
              when "0001" =>
                \$115_n\ := \$v1923\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1922\ := \$arr1644_ptr_take\;
                if \$v1922\(0) = '1' then
                  state_var2258 <= q_wait1921;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1919;
                end if;
              when "0000" =>
                \$116_b\ := \$v1923\(0 to 0);
                \$v1927\ := \$116_b\;
                if \$v1927\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1922\ := \$arr1644_ptr_take\;
                  if \$v1922\(0) = '1' then
                    state_var2258 <= q_wait1921;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1919;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1942 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v176\ := \$arr1644_value\;
              \$v1939\ := \$v176\;
              \$v1940\ := \$v1939\(0 to 3);
              \$v1934\ := \$v1939\(4 to 67);
              case \$v1940\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0011" =>
                \$114_p\ := \$v1934\(0 to 4);
                \$v1936\ := \$114_p\;
                \$v1937\ := \$v1936\(0 to 3);
                \$v1935\ := ""&\$v1936\(4);
                case \$v1937\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0001" =>
                \$115_n\ := \$v1934\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0000" =>
                \$116_b\ := \$v1934\(0 to 0);
                \$v1938\ := \$116_b\;
                if \$v1938\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1958 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v160\ := \$arr1644_value\;
              \$v1955\ := \$v160\;
              \$v1956\ := \$v1955\(0 to 3);
              \$v1950\ := \$v1955\(4 to 67);
              case \$v1956\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                state_var2258 <= \$148_sub572\;
              when "0011" =>
                \$114_p\ := \$v1950\(0 to 4);
                \$v1952\ := \$114_p\;
                \$v1953\ := \$v1952\(0 to 3);
                \$v1951\ := ""&\$v1952\(4);
                case \$v1953\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                state_var2258 <= \$148_sub572\;
              when "0001" =>
                \$115_n\ := \$v1950\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                state_var2258 <= \$148_sub572\;
              when "0000" =>
                \$116_b\ := \$v1950\(0 to 0);
                \$v1954\ := \$116_b\;
                if \$v1954\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_sub572_arg\ := eclat_sub(\$193_n\ & "00000000000000000000000000000001") & debut & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$148_sub572\;
                end if;
              when others =>
                
              end case;
            when pause_getII1969 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v153\ := \$arr1644_value\;
              \$v1966\ := \$v153\;
              \$v1967\ := \$v1966\(0 to 3);
              \$v1961\ := \$v1966\(4 to 67);
              case \$v1967\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1960\ := \$arr1644_ptr_take\;
                if \$v1960\(0) = '1' then
                  state_var2258 <= q_wait1959;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1957;
                end if;
              when "0011" =>
                \$114_p\ := \$v1961\(0 to 4);
                \$v1963\ := \$114_p\;
                \$v1964\ := \$v1963\(0 to 3);
                \$v1962\ := ""&\$v1963\(4);
                case \$v1964\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1960\ := \$arr1644_ptr_take\;
                if \$v1960\(0) = '1' then
                  state_var2258 <= q_wait1959;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1957;
                end if;
              when "0001" =>
                \$115_n\ := \$v1961\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1960\ := \$arr1644_ptr_take\;
                if \$v1960\(0) = '1' then
                  state_var2258 <= q_wait1959;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1957;
                end if;
              when "0000" =>
                \$116_b\ := \$v1961\(0 to 0);
                \$v1965\ := \$116_b\;
                if \$v1965\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1960\ := \$arr1644_ptr_take\;
                  if \$v1960\(0) = '1' then
                    state_var2258 <= q_wait1959;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI1957;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1980 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v150\ := \$arr1644_value\;
              \$v1977\ := \$v150\;
              \$v1978\ := \$v1977\(0 to 3);
              \$v1972\ := \$v1977\(4 to 67);
              case \$v1978\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1971\ := \$arr1644_ptr_take\;
                if \$v1971\(0) = '1' then
                  state_var2258 <= q_wait1970;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1968;
                end if;
              when "0011" =>
                \$114_p\ := \$v1972\(0 to 4);
                \$v1974\ := \$114_p\;
                \$v1975\ := \$v1974\(0 to 3);
                \$v1973\ := ""&\$v1974\(4);
                case \$v1975\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1971\ := \$arr1644_ptr_take\;
                if \$v1971\(0) = '1' then
                  state_var2258 <= q_wait1970;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1968;
                end if;
              when "0001" =>
                \$115_n\ := \$v1972\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1971\ := \$arr1644_ptr_take\;
                if \$v1971\(0) = '1' then
                  state_var2258 <= q_wait1970;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                  state_var2258 <= pause_getI1968;
                end if;
              when "0000" =>
                \$116_b\ := \$v1972\(0 to 0);
                \$v1976\ := \$116_b\;
                if \$v1976\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1971\ := \$arr1644_ptr_take\;
                  if \$v1971\(0) = '1' then
                    state_var2258 <= q_wait1970;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                    state_var2258 <= pause_getI1968;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1987 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v143\ := \$arr1644_value\;
              \$v1984\ := \$v143\;
              \$v1985\ := \$v1984\(0 to 3);
              \$v1983\ := \$v1984\(4 to 67);
              case \$v1985\ is
              when "0001" =>
                a := \$v1983\(0 to 31);
                debut := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1982\ := \$arr1644_ptr_take\;
                if \$v1982\(0) = '1' then
                  state_var2258 <= q_wait1981;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1979;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$121_forever5751634\;
              end case;
            when pause_getII2000 =>
              \$arr1644_ptr_take\(0) := '0';
              \value\ := \$arr1644_value\;
              \$v1997\ := \value\;
              \$v1998\ := \$v1997\(0 to 3);
              \$v1765\ := \$v1997\(4 to 67);
              case \$v1998\ is
              when "0100" =>
                \$v1137\ := \$v1765\(0 to 63);
                \$v1778\ := \$arr1643_ptr_take\;
                if \$v1778\(0) = '1' then
                  state_var2258 <= q_wait1777;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$v1774\ := \$150_vm_run_code547_arg\(32 to 63);
                  \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_add(eclat_add(\$150_vm_run_code547_arg\(160 to 191) & \$193_n\) & "00000000000000000000000000000001") & "00000000000000000000000000000001")));
                  \$arr1643_write_request\ <= '1';
                  \$arr1643_write\ <= "0001" & \$v1774\&X"00000000";
                  state_var2258 <= pause_setI1775;
                end if;
              when "0011" =>
                p := \$v1765\(0 to 4);
                \$v1995\ := p;
                \$v1996\ := \$v1995\(0 to 3);
                \$v1779\ := ""&\$v1995\(4);
                case \$v1996\ is
                when "0101" =>
                  \$v1804\ := eclat_neq(\$193_n\ & "00000000000000000000000000000010");
                  if \$v1804\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2258 <= \$121_forever5751625\;
                  else
                    \$v1803\ := \$arr1644_ptr_take\;
                    if \$v1803\(0) = '1' then
                      state_var2258 <= q_wait1802;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                      state_var2258 <= pause_getI1800;
                    end if;
                  end if;
                when "0110" =>
                  \$v1865\ := eclat_neq(\$193_n\ & "00000000000000000000000000000010");
                  if \$v1865\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2258 <= \$121_forever5751628\;
                  else
                    \$v1864\ := \$arr1644_ptr_take\;
                    if \$v1864\(0) = '1' then
                      state_var2258 <= q_wait1863;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2258 <= pause_getI1861;
                    end if;
                  end if;
                when "0100" =>
                  \$v1884\ := eclat_neq(\$193_n\ & "00000000000000000000000000000010");
                  if \$v1884\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2258 <= \$121_forever5751631\;
                  else
                    \$v1883\ := \$arr1644_ptr_take\;
                    if \$v1883\(0) = '1' then
                      state_var2258 <= q_wait1882;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2258 <= pause_getI1880;
                    end if;
                  end if;
                when "0011" =>
                  \$v1896\ := eclat_lt(\$193_n\ & "00000000000000000000000000000001");
                  if \$v1896\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("pas assez d'arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2258 <= \$121_forever5751633\;
                  else
                    \$v1895\ := \$arr1644_ptr_take\;
                    if \$v1895\(0) = '1' then
                      state_var2258 <= q_wait1894;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                      state_var2258 <= pause_getI1892;
                    end if;
                  end if;
                when "0010" =>
                  \$147_mul571_arg\ := \$193_n\ & "00000000000000000000000000000001" & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$147_mul571\;
                when "0001" =>
                  \$v1990\ := eclat_lt(\$193_n\ & "00000000000000000000000000000010");
                  if \$v1990\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut 2 arguments pour la soustraction"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2258 <= \$121_forever5751635\;
                  else
                    \$v1989\ := \$arr1644_ptr_take\;
                    if \$v1989\(0) = '1' then
                      state_var2258 <= q_wait1988;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                      state_var2258 <= pause_getI1986;
                    end if;
                  end if;
                when "0000" =>
                  \$149_add573_arg\ := \$193_n\ & "00000000000000000000000000000000" & \$150_vm_run_code547_arg\(0 to 31);
                  state_var2258 <= \$149_add573\;
                when others =>
                  \$166\ := \$150_vm_run_code547_arg\(0 to 293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                end case;
              when others =>
                \$166\ := \$150_vm_run_code547_arg\(0 to 293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              end case;
            when pause_getII2013 =>
              \$arr1647_ptr_take\(0) := '0';
              \$v1476\ := \$arr1647_value\;
              \$v2011\ := \$arr1644_ptr_take\;
              if \$v2011\(0) = '1' then
                state_var2258 <= q_wait2010;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$v1476\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= v;
                state_var2258 <= pause_setI2008;
              end if;
            when pause_getII2017 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2015\ := \$arr1647_ptr_take\;
              if \$v2015\(0) = '1' then
                state_var2258 <= q_wait2014;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2012;
              end if;
            when pause_getII2024 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2021\ := v;
              \$v2022\ := \$v2021\(0 to 3);
              \$v2020\ := \$v2021\(4 to 67);
              case \$v2022\ is
              when "0000" =>
                x := \$v2020\(0 to 0);
                condition := x;
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & 
                eclat_if(condition & \$150_vm_run_code547_arg\(64 to 95) & eclat_sub(\$196_l\ & "00000000000000000000000000000001")) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when others =>
                condition := eclat_false;
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & 
                eclat_if(condition & \$150_vm_run_code547_arg\(64 to 95) & eclat_sub(\$196_l\ & "00000000000000000000000000000001")) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              end case;
            when pause_getII2031 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2028\ := v;
              \$v2029\ := \$v2028\(0 to 3);
              \$v2027\ := \$v2028\(4 to 67);
              case \$v2029\ is
              when "0000" =>
                x := \$v2027\(0 to 0);
                cond := x;
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$197_l\ & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(64 to 95)) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when others =>
                cond := eclat_false;
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$197_l\ & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(64 to 95)) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              end case;
            when pause_getII2039 =>
              \$arr1644_ptr_take\(0) := '0';
              var := \$arr1644_value\;
              \$v2037\ := \$arr1643_ptr_take\;
              if \$v2037\(0) = '1' then
                state_var2258 <= q_wait2036;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$198_i\)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= var;
                state_var2258 <= pause_setI2034;
              end if;
            when pause_getII2047 =>
              \$arr1643_ptr_take\(0) := '0';
              local_value := \$arr1643_value\;
              \$v2045\ := \$arr1644_ptr_take\;
              if \$v2045\(0) = '1' then
                state_var2258 <= q_wait2044;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= local_value;
                state_var2258 <= pause_setI2042;
              end if;
            when pause_getII2058 =>
              \$arr1643_ptr_take\(0) := '0';
              \$v213\ := \$arr1643_value\;
              \$v2055\ := \$v213\;
              \$v2056\ := \$v2055\(0 to 3);
              \$v2050\ := \$v2055\(4 to 67);
              case \$v2056\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2258 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                  state_var2258 <= pause_getI2046;
                end if;
              when "0011" =>
                \$114_p\ := \$v2050\(0 to 4);
                \$v2052\ := \$114_p\;
                \$v2053\ := \$v2052\(0 to 3);
                \$v2051\ := ""&\$v2052\(4);
                case \$v2053\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2258 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                  state_var2258 <= pause_getI2046;
                end if;
              when "0001" =>
                \$115_n\ := \$v2050\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2258 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                  state_var2258 <= pause_getI2046;
                end if;
              when "0000" =>
                \$116_b\ := \$v2050\(0 to 0);
                \$v2054\ := \$116_b\;
                if \$v2054\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2258 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                    state_var2258 <= pause_getI2046;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2066 =>
              \$arr1645_ptr_take\(0) := '0';
              \$v217\ := \$arr1645_value\;
              \$v2064\ := \$arr1644_ptr_take\;
              if \$v2064\(0) = '1' then
                state_var2258 <= q_wait2063;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$v217\;
                state_var2258 <= pause_setI2061;
              end if;
            when pause_getII2074 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v221\ := \$arr1644_value\;
              \$v2072\ := \$arr1645_ptr_take\;
              if \$v2072\(0) = '1' then
                state_var2258 <= q_wait2071;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr_write\ <= to_integer(unsigned(\$202_i\));
                \$arr1645_write_request\ <= '1';
                \$arr1645_write\ <= \$v221\;
                state_var2258 <= pause_setI2069;
              end if;
            when pause_getII2085 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v229\ := \$arr1644_value\;
              \$v2082\ := \$v229\;
              \$v2083\ := \$v2082\(0 to 3);
              \$v2077\ := \$v2082\(4 to 67);
              case \$v2083\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0011" =>
                \$114_p\ := \$v2077\(0 to 4);
                \$v2079\ := \$114_p\;
                \$v2080\ := \$v2079\(0 to 3);
                \$v2078\ := ""&\$v2079\(4);
                case \$v2080\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0001" =>
                \$115_n\ := \$v2077\(0 to 31);
                eclat_print_int(\$115_n\);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0000" =>
                \$116_b\ := \$v2077\(0 to 0);
                \$v2081\ := \$116_b\;
                if \$v2081\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & eclat_true;
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2096 =>
              \$arr1646_ptr_take\(0) := '0';
              \$192_instr\ := \$arr1646_value\;
              \$v2093\ := \$192_instr\;
              \$v2094\ := \$v2093\(0 to 3);
              \$v1764\ := \$v2093\(4 to 71);
              case \$v2094\ is
              when "1000" =>
                \$193_n\ := \$v1764\(0 to 31);
                \$v2002\ := \$arr1644_ptr_take\;
                if \$v2002\(0) = '1' then
                  state_var2258 <= q_wait2001;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI1999;
                end if;
              when "0110" =>
                \$194_l\ := \$v1764\(0 to 31);
                \$v2007\ := \$arr1644_ptr_take\;
                if \$v2007\(0) = '1' then
                  state_var2258 <= q_wait2006;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v2003\ := \$194_l\ & \$150_vm_run_code547_arg\(32 to 63);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0100" & \$v2003\;
                  state_var2258 <= pause_setI2004;
                end if;
              when "1001" =>
                \$v2019\ := \$arr1644_ptr_take\;
                if \$v2019\(0) = '1' then
                  state_var2258 <= q_wait2018;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI2016;
                end if;
              when "1100" =>
                \$196_l\ := \$v1764\(0 to 31);
                \$v2026\ := \$arr1644_ptr_take\;
                if \$v2026\(0) = '1' then
                  state_var2258 <= q_wait2025;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI2023;
                end if;
              when "1011" =>
                \$197_l\ := \$v1764\(0 to 31);
                \$v2033\ := \$arr1644_ptr_take\;
                if \$v2033\(0) = '1' then
                  state_var2258 <= q_wait2032;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI2030;
                end if;
              when "0011" =>
                \$198_i\ := \$v1764\(0 to 31);
                \$v2041\ := \$arr1644_ptr_take\;
                if \$v2041\(0) = '1' then
                  state_var2258 <= q_wait2040;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI2038;
                end if;
              when "1010" =>
                \$199_l\ := \$v1764\(0 to 31);
                \$166\ := \$150_vm_run_code547_arg\(0 to 31) & \$150_vm_run_code547_arg\(32 to 63) & eclat_sub(\$199_l\ & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0100" =>
                \$200_i\ := \$v1764\(0 to 31);
                eclat_print_string(of_string("env "));
                
                eclat_print_int(\$150_vm_run_code547_arg\(32 to 63));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2060\ := \$arr1643_ptr_take\;
                if \$v2060\(0) = '1' then
                  state_var2258 <= q_wait2059;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                  state_var2258 <= pause_getI2057;
                end if;
              when "0010" =>
                \$201_i\ := \$v1764\(0 to 31);
                \$v2068\ := \$arr1645_ptr_take\;
                if \$v2068\(0) = '1' then
                  state_var2258 <= q_wait2067;
                else
                  \$arr1645_ptr_take\(0) := '1';
                  \$arr1645_ptr\ <= to_integer(unsigned(\$201_i\));
                  state_var2258 <= pause_getI2065;
                end if;
              when "0001" =>
                \$202_i\ := \$v1764\(0 to 31);
                \$v2076\ := \$arr1644_ptr_take\;
                if \$v2076\(0) = '1' then
                  state_var2258 <= q_wait2075;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2258 <= pause_getI2073;
                end if;
              when "0000" =>
                \$166\ := \$150_vm_run_code547_arg\(0 to 31) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & eclat_add(\$150_vm_run_code547_arg\(128 to 159) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0111" =>
                \$v2088\ := eclat_eq(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & "00000000000000000000000000000000");
                if \$v2088\(0) = '1' then
                  \$v2087\ := \$arr1644_ptr_take\;
                  if \$v2087\(0) = '1' then
                    state_var2258 <= q_wait2086;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2258 <= pause_getI2084;
                  end if;
                else
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                end if;
              when "0101" =>
                \$205_v\ := \$v1764\(0 to 67);
                \$v2092\ := \$arr1644_ptr_take\;
                if \$v2092\(0) = '1' then
                  state_var2258 <= q_wait2091;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= \$205_v\;
                  state_var2258 <= pause_setI2089;
                end if;
              when others =>
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2258 <= \$209_forever5741620\;
              end case;
            when pause_setI1720 =>
              \$arr1643_write_request\ <= '0';
              state_var2258 <= pause_setII1721;
            when pause_setI1766 =>
              \$arr1647_write_request\ <= '0';
              state_var2258 <= pause_setII1767;
            when pause_setI1770 =>
              \$arr1647_write_request\ <= '0';
              state_var2258 <= pause_setII1771;
            when pause_setI1775 =>
              \$arr1643_write_request\ <= '0';
              state_var2258 <= pause_setII1776;
            when pause_setI1780 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1781;
            when pause_setI1814 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1815;
            when pause_setI1866 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1867;
            when pause_setI1885 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1886;
            when pause_setI1897 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1898;
            when pause_setI1946 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1947;
            when pause_setI1991 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII1992;
            when pause_setI2004 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII2005;
            when pause_setI2008 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII2009;
            when pause_setI2034 =>
              \$arr1643_write_request\ <= '0';
              state_var2258 <= pause_setII2035;
            when pause_setI2042 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII2043;
            when pause_setI2061 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII2062;
            when pause_setI2069 =>
              \$arr1645_write_request\ <= '0';
              state_var2258 <= pause_setII2070;
            when pause_setI2089 =>
              \$arr1644_write_request\ <= '0';
              state_var2258 <= pause_setII2090;
            when pause_setII1721 =>
              \$arr1643_ptr_take\(0) := '0';
              eclat_print_string(of_string("copy heap["));
              
              eclat_print_int(\$144_copy_args_to_heap544_arg\(64 to 95));
              
              eclat_print_string(of_string("] <-"));
              
              \$v1719\ := \$arr1644_ptr_take\;
              if \$v1719\(0) = '1' then
                state_var2258 <= q_wait1718;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$144_copy_args_to_heap544_arg\(32 to 63) & \$144_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1716;
              end if;
            when pause_setII1767 =>
              \$arr1647_ptr_take\(0) := '0';
              \$166\ := eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(160 to 191) & eclat_sub(\$v1137\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$150_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(128 to 159) & eclat_add(eclat_add(\$150_vm_run_code547_arg\(160 to 191) & \$193_n\) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII1771 =>
              \$arr1647_ptr_take\(0) := '0';
              \$v1769\ := \$arr1647_ptr_take\;
              if \$v1769\(0) = '1' then
                state_var2258 <= q_wait1768;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001") & \$v1137\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127);
                state_var2258 <= pause_setI1766;
              end if;
            when pause_setII1776 =>
              \$arr1643_ptr_take\(0) := '0';
              \$144_copy_args_to_heap544_arg\ := \$193_n\ & \$150_vm_run_code547_arg\(0 to 31) & \$150_vm_run_code547_arg\(160 to 191);
              state_var2258 <= \$144_copy_args_to_heap544\;
            when pause_setII1781 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII1815 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_string(of_string("ICIIIIIIIII"));
              
              \$v1812\ := eclat_gt(fst_operand & scd_operand);
              \$v1810\ := "0000" & \$v1812\&"000"& X"000000000000000";
              \$v1811\ := \$v1810\(0 to 3);
              \$v1805\ := \$v1810\(4 to 67);
              case \$v1811\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0011" =>
                \$114_p\ := \$v1805\(0 to 4);
                \$v1807\ := \$114_p\;
                \$v1808\ := \$v1807\(0 to 3);
                \$v1806\ := ""&\$v1807\(4);
                case \$v1808\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0001" =>
                \$115_n\ := \$v1805\(0 to 31);
                eclat_print_int(\$115_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                \$v1763\ := ""&\$166\(293);
                if \$v1763\(0) = '1' then
                  \$150_vm_run_code547_result\ := eclat_unit;
                  result1706 := \$150_vm_run_code547_result\;
                  rdy1707 := eclat_true;
                  state_var2258 <= compute1708;
                else
                  \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                  state_var2258 <= \$150_vm_run_code547\;
                end if;
              when "0000" =>
                \$116_b\ := \$v1805\(0 to 0);
                \$v1809\ := \$116_b\;
                if \$v1809\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
                  \$v1763\ := ""&\$166\(293);
                  if \$v1763\(0) = '1' then
                    \$150_vm_run_code547_result\ := eclat_unit;
                    result1706 := \$150_vm_run_code547_result\;
                    rdy1707 := eclat_true;
                    state_var2258 <= compute1708;
                  else
                    \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                    state_var2258 <= \$150_vm_run_code547\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_setII1867 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII1886 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII1898 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII1947 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_string(of_string("le resultat :stack["));
              
              eclat_print_int(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001"));
              
              eclat_print_string(of_string("] <-"));
              
              \$v1944\ := \$arr1644_ptr_take\;
              if \$v1944\(0) = '1' then
                state_var2258 <= q_wait1943;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1941;
              end if;
            when pause_setII1992 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2005 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_add(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2009 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_add(\$v1476\(0 to 31) & "00000000000000000000000000000001") & \$v1476\(32 to 63) & \$v1476\(64 to 95) & \$v1476\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2035 =>
              \$arr1643_ptr_take\(0) := '0';
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2043 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_add(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2062 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_add(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2070 =>
              \$arr1645_ptr_take\(0) := '0';
              \$166\ := eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when pause_setII2090 =>
              \$arr1644_ptr_take\(0) := '0';
              \$166\ := eclat_add(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127) & \$150_vm_run_code547_arg\(128 to 159) & \$150_vm_run_code547_arg\(160 to 191) & \$150_vm_run_code547_arg\(192 to 292) & ""&\$150_vm_run_code547_arg\(293);
              \$v1763\ := ""&\$166\(293);
              if \$v1763\(0) = '1' then
                \$150_vm_run_code547_result\ := eclat_unit;
                result1706 := \$150_vm_run_code547_result\;
                rdy1707 := eclat_true;
                state_var2258 <= compute1708;
              else
                \$150_vm_run_code547_arg\ := \$166\(0 to 31) & \$166\(32 to 63) & eclat_add(\$166\(64 to 95) & "00000000000000000000000000000001") & \$166\(96 to 127) & \$166\(128 to 159) & \$166\(160 to 191) & \$166\(192 to 292) & ""&\$166\(293) & ""&\$150_vm_run_code547_arg\(294);
                state_var2258 <= \$150_vm_run_code547\;
              end if;
            when q_wait1718 =>
              \$v1719\ := \$arr1644_ptr_take\;
              if \$v1719\(0) = '1' then
                state_var2258 <= q_wait1718;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$144_copy_args_to_heap544_arg\(32 to 63) & \$144_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1716;
              end if;
            when q_wait1722 =>
              \$v1723\ := \$arr1643_ptr_take\;
              if \$v1723\(0) = '1' then
                state_var2258 <= q_wait1722;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(\$144_copy_args_to_heap544_arg\(64 to 95)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= \$404\;
                state_var2258 <= pause_setI1720;
              end if;
            when q_wait1726 =>
              \$v1727\ := \$arr1644_ptr_take\;
              if \$v1727\(0) = '1' then
                state_var2258 <= q_wait1726;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$144_copy_args_to_heap544_arg\(32 to 63) & \$144_copy_args_to_heap544_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1724;
              end if;
            when q_wait1736 =>
              \$v1737\ := \$arr1644_ptr_take\;
              if \$v1737\(0) = '1' then
                state_var2258 <= q_wait1736;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_div570_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_div570_arg\(0 to 31))));
                state_var2258 <= pause_getI1734;
              end if;
            when q_wait1744 =>
              \$v1745\ := \$arr1644_ptr_take\;
              if \$v1745\(0) = '1' then
                state_var2258 <= q_wait1744;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_mul571_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_mul571_arg\(0 to 31))));
                state_var2258 <= pause_getI1742;
              end if;
            when q_wait1752 =>
              \$v1753\ := \$arr1644_ptr_take\;
              if \$v1753\(0) = '1' then
                state_var2258 <= q_wait1752;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_sub572_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_sub572_arg\(0 to 31))));
                state_var2258 <= pause_getI1750;
              end if;
            when q_wait1760 =>
              \$v1761\ := \$arr1644_ptr_take\;
              if \$v1761\(0) = '1' then
                state_var2258 <= q_wait1760;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_add573_arg\(64 to 95) & "00000000000000000000000000000001") & \$149_add573_arg\(0 to 31))));
                state_var2258 <= pause_getI1758;
              end if;
            when q_wait1768 =>
              \$v1769\ := \$arr1647_ptr_take\;
              if \$v1769\(0) = '1' then
                state_var2258 <= q_wait1768;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001") & \$v1137\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127);
                state_var2258 <= pause_setI1766;
              end if;
            when q_wait1772 =>
              \$v1773\ := \$arr1647_ptr_take\;
              if \$v1773\(0) = '1' then
                state_var2258 <= q_wait1772;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(96 to 127)));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001") & \$150_vm_run_code547_arg\(32 to 63) & \$150_vm_run_code547_arg\(64 to 95) & \$150_vm_run_code547_arg\(96 to 127);
                state_var2258 <= pause_setI1770;
              end if;
            when q_wait1777 =>
              \$v1778\ := \$arr1643_ptr_take\;
              if \$v1778\(0) = '1' then
                state_var2258 <= q_wait1777;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$v1774\ := \$150_vm_run_code547_arg\(32 to 63);
                \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_add(eclat_add(\$150_vm_run_code547_arg\(160 to 191) & \$193_n\) & "00000000000000000000000000000001") & "00000000000000000000000000000001")));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= "0001" & \$v1774\&X"00000000";
                state_var2258 <= pause_setI1775;
              end if;
            when q_wait1782 =>
              \$v1783\ := \$arr1644_ptr_take\;
              if \$v1783\(0) = '1' then
                state_var2258 <= q_wait1782;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001") & \$193_n\)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                state_var2258 <= pause_setI1780;
              end if;
            when q_wait1798 =>
              \$v1799\ := \$arr1644_ptr_take\;
              if \$v1799\(0) = '1' then
                state_var2258 <= q_wait1798;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2258 <= pause_getI1796;
              end if;
            when q_wait1802 =>
              \$v1803\ := \$arr1644_ptr_take\;
              if \$v1803\(0) = '1' then
                state_var2258 <= q_wait1802;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2258 <= pause_getI1800;
              end if;
            when q_wait1816 =>
              \$v1817\ := \$arr1644_ptr_take\;
              if \$v1817\(0) = '1' then
                state_var2258 <= q_wait1816;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v1813\ := eclat_gt(fst_operand & scd_operand);
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0000" & \$v1813\&"000"& X"000000000000000";
                state_var2258 <= pause_setI1814;
              end if;
            when q_wait1827 =>
              \$v1828\ := \$arr1644_ptr_take\;
              if \$v1828\(0) = '1' then
                state_var2258 <= q_wait1827;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1825;
              end if;
            when q_wait1838 =>
              \$v1839\ := \$arr1644_ptr_take\;
              if \$v1839\(0) = '1' then
                state_var2258 <= q_wait1838;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2258 <= pause_getI1836;
              end if;
            when q_wait1849 =>
              \$v1850\ := \$arr1644_ptr_take\;
              if \$v1850\(0) = '1' then
                state_var2258 <= q_wait1849;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2258 <= pause_getI1847;
              end if;
            when q_wait1856 =>
              \$v1857\ := \$arr1644_ptr_take\;
              if \$v1857\(0) = '1' then
                state_var2258 <= q_wait1856;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2258 <= pause_getI1854;
              end if;
            when q_wait1863 =>
              \$v1864\ := \$arr1644_ptr_take\;
              if \$v1864\(0) = '1' then
                state_var2258 <= q_wait1863;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2258 <= pause_getI1861;
              end if;
            when q_wait1868 =>
              \$v1869\ := \$arr1644_ptr_take\;
              if \$v1869\(0) = '1' then
                state_var2258 <= q_wait1868;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2258 <= pause_setI1866;
              end if;
            when q_wait1875 =>
              \$v1876\ := \$arr1644_ptr_take\;
              if \$v1876\(0) = '1' then
                state_var2258 <= q_wait1875;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2258 <= pause_getI1873;
              end if;
            when q_wait1882 =>
              \$v1883\ := \$arr1644_ptr_take\;
              if \$v1883\(0) = '1' then
                state_var2258 <= q_wait1882;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2258 <= pause_getI1880;
              end if;
            when q_wait1887 =>
              \$v1888\ := \$arr1644_ptr_take\;
              if \$v1888\(0) = '1' then
                state_var2258 <= q_wait1887;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2258 <= pause_setI1885;
              end if;
            when q_wait1894 =>
              \$v1895\ := \$arr1644_ptr_take\;
              if \$v1895\(0) = '1' then
                state_var2258 <= q_wait1894;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1892;
              end if;
            when q_wait1899 =>
              \$v1900\ := \$arr1644_ptr_take\;
              if \$v1900\(0) = '1' then
                state_var2258 <= q_wait1899;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2258 <= pause_setI1897;
              end if;
            when q_wait1910 =>
              \$v1911\ := \$arr1644_ptr_take\;
              if \$v1911\(0) = '1' then
                state_var2258 <= q_wait1910;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1908;
              end if;
            when q_wait1921 =>
              \$v1922\ := \$arr1644_ptr_take\;
              if \$v1922\(0) = '1' then
                state_var2258 <= q_wait1921;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                state_var2258 <= pause_getI1919;
              end if;
            when q_wait1932 =>
              \$v1933\ := \$arr1644_ptr_take\;
              if \$v1933\(0) = '1' then
                state_var2258 <= q_wait1932;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1930;
              end if;
            when q_wait1943 =>
              \$v1944\ := \$arr1644_ptr_take\;
              if \$v1944\(0) = '1' then
                state_var2258 <= q_wait1943;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1941;
              end if;
            when q_wait1948 =>
              \$v1949\ := \$arr1644_ptr_take\;
              if \$v1949\(0) = '1' then
                state_var2258 <= q_wait1948;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v1945\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & \$v1945\&X"00000000";
                state_var2258 <= pause_setI1946;
              end if;
            when q_wait1959 =>
              \$v1960\ := \$arr1644_ptr_take\;
              if \$v1960\(0) = '1' then
                state_var2258 <= q_wait1959;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1957;
              end if;
            when q_wait1970 =>
              \$v1971\ := \$arr1644_ptr_take\;
              if \$v1971\(0) = '1' then
                state_var2258 <= q_wait1970;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\)));
                state_var2258 <= pause_getI1968;
              end if;
            when q_wait1981 =>
              \$v1982\ := \$arr1644_ptr_take\;
              if \$v1982\(0) = '1' then
                state_var2258 <= q_wait1981;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1979;
              end if;
            when q_wait1988 =>
              \$v1989\ := \$arr1644_ptr_take\;
              if \$v1989\(0) = '1' then
                state_var2258 <= q_wait1988;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1986;
              end if;
            when q_wait1993 =>
              \$v1994\ := \$arr1644_ptr_take\;
              if \$v1994\(0) = '1' then
                state_var2258 <= q_wait1993;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & \$193_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2258 <= pause_setI1991;
              end if;
            when q_wait2001 =>
              \$v2002\ := \$arr1644_ptr_take\;
              if \$v2002\(0) = '1' then
                state_var2258 <= q_wait2001;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI1999;
              end if;
            when q_wait2006 =>
              \$v2007\ := \$arr1644_ptr_take\;
              if \$v2007\(0) = '1' then
                state_var2258 <= q_wait2006;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v2003\ := \$194_l\ & \$150_vm_run_code547_arg\(32 to 63);
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0100" & \$v2003\;
                state_var2258 <= pause_setI2004;
              end if;
            when q_wait2010 =>
              \$v2011\ := \$arr1644_ptr_take\;
              if \$v2011\(0) = '1' then
                state_var2258 <= q_wait2010;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$v1476\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= v;
                state_var2258 <= pause_setI2008;
              end if;
            when q_wait2014 =>
              \$v2015\ := \$arr1647_ptr_take\;
              if \$v2015\(0) = '1' then
                state_var2258 <= q_wait2014;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(96 to 127) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2012;
              end if;
            when q_wait2018 =>
              \$v2019\ := \$arr1644_ptr_take\;
              if \$v2019\(0) = '1' then
                state_var2258 <= q_wait2018;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2016;
              end if;
            when q_wait2025 =>
              \$v2026\ := \$arr1644_ptr_take\;
              if \$v2026\(0) = '1' then
                state_var2258 <= q_wait2025;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2023;
              end if;
            when q_wait2032 =>
              \$v2033\ := \$arr1644_ptr_take\;
              if \$v2033\(0) = '1' then
                state_var2258 <= q_wait2032;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2030;
              end if;
            when q_wait2036 =>
              \$v2037\ := \$arr1643_ptr_take\;
              if \$v2037\(0) = '1' then
                state_var2258 <= q_wait2036;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$198_i\)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= var;
                state_var2258 <= pause_setI2034;
              end if;
            when q_wait2040 =>
              \$v2041\ := \$arr1644_ptr_take\;
              if \$v2041\(0) = '1' then
                state_var2258 <= q_wait2040;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2038;
              end if;
            when q_wait2044 =>
              \$v2045\ := \$arr1644_ptr_take\;
              if \$v2045\(0) = '1' then
                state_var2258 <= q_wait2044;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= local_value;
                state_var2258 <= pause_setI2042;
              end if;
            when q_wait2048 =>
              \$v2049\ := \$arr1643_ptr_take\;
              if \$v2049\(0) = '1' then
                state_var2258 <= q_wait2048;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                state_var2258 <= pause_getI2046;
              end if;
            when q_wait2059 =>
              \$v2060\ := \$arr1643_ptr_take\;
              if \$v2060\(0) = '1' then
                state_var2258 <= q_wait2059;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$150_vm_run_code547_arg\(32 to 63) & \$200_i\)));
                state_var2258 <= pause_getI2057;
              end if;
            when q_wait2063 =>
              \$v2064\ := \$arr1644_ptr_take\;
              if \$v2064\(0) = '1' then
                state_var2258 <= q_wait2063;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$v217\;
                state_var2258 <= pause_setI2061;
              end if;
            when q_wait2067 =>
              \$v2068\ := \$arr1645_ptr_take\;
              if \$v2068\(0) = '1' then
                state_var2258 <= q_wait2067;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr\ <= to_integer(unsigned(\$201_i\));
                state_var2258 <= pause_getI2065;
              end if;
            when q_wait2071 =>
              \$v2072\ := \$arr1645_ptr_take\;
              if \$v2072\(0) = '1' then
                state_var2258 <= q_wait2071;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr_write\ <= to_integer(unsigned(\$202_i\));
                \$arr1645_write_request\ <= '1';
                \$arr1645_write\ <= \$v221\;
                state_var2258 <= pause_setI2069;
              end if;
            when q_wait2075 =>
              \$v2076\ := \$arr1644_ptr_take\;
              if \$v2076\(0) = '1' then
                state_var2258 <= q_wait2075;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2073;
              end if;
            when q_wait2086 =>
              \$v2087\ := \$arr1644_ptr_take\;
              if \$v2087\(0) = '1' then
                state_var2258 <= q_wait2086;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$150_vm_run_code547_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2258 <= pause_getI2084;
              end if;
            when q_wait2091 =>
              \$v2092\ := \$arr1644_ptr_take\;
              if \$v2092\(0) = '1' then
                state_var2258 <= q_wait2091;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$205_v\;
                state_var2258 <= pause_setI2089;
              end if;
            when q_wait2097 =>
              \$v2098\ := \$arr1646_ptr_take\;
              if \$v2098\(0) = '1' then
                state_var2258 <= q_wait2097;
              else
                \$arr1646_ptr_take\(0) := '1';
                \$arr1646_ptr\ <= to_integer(unsigned(\$150_vm_run_code547_arg\(64 to 95)));
                state_var2258 <= pause_getI2095;
              end if;
            when compute1708 =>
              rdy1707 := eclat_false;
              eclat_print_string(of_string("START (cy="));
              
              eclat_print_int(\$136_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              \$v2100\ := eclat_unit;
              \$150_vm_run_code547_arg\ := "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & eclat_false & "00000000000000000000000000000000" & "0010" & \$v2100\&"000"& X"000000000000000" & eclat_false & argument;
              state_var2258 <= \$150_vm_run_code547\;
            end case;
            \$v2102\ := eclat_not(rdy1707);
            if \$v2102\(0) = '1' then
              result1706 := eclat_unit;
            end if;
            \$137\ := result1706 & rdy1707;
            \$v1705\ := ""&\$137\(1);
            if \$v1705\(0) = '1' then
              eclat_print_string(of_string("END (cy="));
              
              eclat_print_int(\$136_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              result1648 := eclat_unit;
              eclat_print_newline(eclat_unit);
              
              rdy1649 := eclat_true;
              \state\ <= compute1650;
            else
              result1648 := eclat_unit;
              rdy1649 := eclat_true;
              \state\ <= compute1650;
            end if;
          end case;
          
          result <= result1648;
          rdy <= rdy1649;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
