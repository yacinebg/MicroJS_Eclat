-- code generated from the following source code:
--   ../vm/fail.ecl
--   ../vm/value.ecl
--   ../vm/ram.ecl
--   ../vm/frames.ecl
--   ../vm/vm.ecl
--   ../vm/main.ecl
--
-- with the following command:
--
--    ./eclat -arg=true -relax -notyB ../vm/fail.ecl ../vm/value.ecl ../vm/ram.ecl ../vm/frames.ecl ../vm/vm.ecl ../vm/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute1650, \$127_copy_args_to_heap518\, \$128_pow542\, \$129_div543\, \$130_mul544\, \$131_sub545\, \$132_add546\, \$615_forever5481612\, \$640_forever5481611\, \$665_forever5481610\, \$689_forever5481608\, \$698_forever5481609\, pause_getI1655, pause_getI1665, pause_getI1673, pause_getI1681, pause_getI1689, pause_getII1656, pause_getII1666, pause_getII1674, pause_getII1682, pause_getII1690, pause_setI1651, pause_setII1652, q_wait1653, q_wait1657, q_wait1667, q_wait1675, q_wait1683, q_wait1691);
  signal \state\: t_state;
  type t_state_var2250 is (compute2113, \$400_copy_args_to_heap518\, \$401_pow542\, \$402_div543\, \$403_mul544\, \$404_sub545\, \$405_add546\, \$462_forever5481642\, \$466_forever5481636\, \$491_forever5481641\, \$495_forever5481636\, \$520_forever5481640\, \$524_forever5481636\, \$548_forever5481638\, \$552_forever5481636\, \$561_forever5481639\, \$565_forever5481636\, pause_getI2118, pause_getI2128, pause_getI2136, pause_getI2144, pause_getI2152, pause_getII2119, pause_getII2129, pause_getII2137, pause_getII2145, pause_getII2153, pause_setI2114, pause_setI2158, pause_setI2163, pause_setI2168, pause_setI2174, pause_setI2180, pause_setI2185, pause_setI2190, pause_setI2195, pause_setI2201, pause_setI2206, pause_setI2211, pause_setI2218, pause_setI2223, pause_setI2228, pause_setI2233, pause_setI2238, pause_setII2115, pause_setII2159, pause_setII2164, pause_setII2169, pause_setII2175, pause_setII2181, pause_setII2186, pause_setII2191, pause_setII2196, pause_setII2202, pause_setII2207, pause_setII2212, pause_setII2219, pause_setII2224, pause_setII2229, pause_setII2234, pause_setII2239, q_wait2116, q_wait2120, q_wait2130, q_wait2138, q_wait2146, q_wait2154, q_wait2160, q_wait2165, q_wait2170, q_wait2176, q_wait2182, q_wait2187, q_wait2192, q_wait2197, q_wait2203, q_wait2208, q_wait2213, q_wait2220, q_wait2225, q_wait2230, q_wait2235, q_wait2240);
  signal state_var2250: t_state_var2250;
  type t_state_var2249 is (compute2110);
  signal state_var2249: t_state_var2249;
  type t_state_var2248 is (compute2105);
  signal state_var2248: t_state_var2248;
  type t_state_var2247 is (compute1697, \$117_forever5471614\, \$117_forever5471621\, \$117_forever5471622\, \$117_forever5471623\, \$117_forever5471624\, \$120_forever5481613\, \$120_forever5481625\, \$120_forever5481626\, \$120_forever5481627\, \$120_forever5481628\, \$120_forever5481629\, \$120_forever5481630\, \$120_forever5481631\, \$120_forever5481632\, \$120_forever5481633\, \$120_forever5481634\, \$120_forever5481635\, \$143_copy_args_to_heap518\, \$144_pow542\, \$145_div543\, \$146_mul544\, \$147_sub545\, \$148_add546\, \$149_vm_run_code521\, \$208_forever5471620\, \$212_forever5471614\, \$258_forever5481619\, \$262_forever5481613\, \$287_forever5481618\, \$291_forever5481613\, \$316_forever5481617\, \$320_forever5481613\, \$344_forever5481615\, \$348_forever5481613\, \$357_forever5481616\, \$361_forever5481613\, pause_getI1702, pause_getI1712, pause_getI1720, pause_getI1728, pause_getI1736, pause_getI1774, pause_getI1778, pause_getI1803, pause_getI1814, pause_getI1825, pause_getI1832, pause_getI1839, pause_getI1851, pause_getI1858, pause_getI1870, pause_getI1886, pause_getI1897, pause_getI1908, pause_getI1924, pause_getI1935, pause_getI1946, pause_getI1953, pause_getI1969, pause_getI1980, pause_getI1991, pause_getI1999, pause_getI2012, pause_getI2016, pause_getI2023, pause_getI2030, pause_getI2038, pause_getI2046, pause_getI2057, pause_getI2065, pause_getI2073, pause_getI2084, pause_getI2095, pause_getII1703, pause_getII1713, pause_getII1721, pause_getII1729, pause_getII1737, pause_getII1775, pause_getII1779, pause_getII1804, pause_getII1815, pause_getII1826, pause_getII1833, pause_getII1840, pause_getII1852, pause_getII1859, pause_getII1871, pause_getII1887, pause_getII1898, pause_getII1909, pause_getII1925, pause_getII1936, pause_getII1947, pause_getII1954, pause_getII1970, pause_getII1981, pause_getII1992, pause_getII2000, pause_getII2013, pause_getII2017, pause_getII2024, pause_getII2031, pause_getII2039, pause_getII2047, pause_getII2058, pause_getII2066, pause_getII2074, pause_getII2085, pause_getII2096, pause_setI1698, pause_setI1744, pause_setI1748, pause_setI1753, pause_setI1758, pause_setI1792, pause_setI1844, pause_setI1863, pause_setI1875, pause_setI1913, pause_setI1958, pause_setI2004, pause_setI2008, pause_setI2034, pause_setI2042, pause_setI2061, pause_setI2069, pause_setI2089, pause_setII1699, pause_setII1745, pause_setII1749, pause_setII1754, pause_setII1759, pause_setII1793, pause_setII1845, pause_setII1864, pause_setII1876, pause_setII1914, pause_setII1959, pause_setII2005, pause_setII2009, pause_setII2035, pause_setII2043, pause_setII2062, pause_setII2070, pause_setII2090, q_wait1700, q_wait1704, q_wait1714, q_wait1722, q_wait1730, q_wait1738, q_wait1746, q_wait1750, q_wait1755, q_wait1760, q_wait1776, q_wait1780, q_wait1794, q_wait1805, q_wait1816, q_wait1827, q_wait1834, q_wait1841, q_wait1846, q_wait1853, q_wait1860, q_wait1865, q_wait1872, q_wait1877, q_wait1888, q_wait1899, q_wait1910, q_wait1915, q_wait1926, q_wait1937, q_wait1948, q_wait1955, q_wait1960, q_wait1971, q_wait1982, q_wait1993, q_wait2001, q_wait2006, q_wait2010, q_wait2014, q_wait2018, q_wait2025, q_wait2032, q_wait2036, q_wait2040, q_wait2044, q_wait2048, q_wait2059, q_wait2063, q_wait2067, q_wait2071, q_wait2075, q_wait2086, q_wait2091, q_wait2097);
  signal state_var2247: t_state_var2247;
  type array_value_68 is array (natural range <>) of value(0 to 67);
  type array_value_72 is array (natural range <>) of value(0 to 71);
  type array_value_128 is array (natural range <>) of value(0 to 127);
  signal arr1643 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1643_value\ : value(0 to 67);
  signal \$arr1643_ptr\ : natural range 0 to 99;
  signal \$arr1643_ptr_write\ : natural range 0 to 99;
  signal \$arr1643_write\ : value(0 to 67);
  signal \$arr1643_write_request\ : std_logic := '0';
  signal arr1644 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1644_value\ : value(0 to 67);
  signal \$arr1644_ptr\ : natural range 0 to 99;
  signal \$arr1644_ptr_write\ : natural range 0 to 99;
  signal \$arr1644_write\ : value(0 to 67);
  signal \$arr1644_write_request\ : std_logic := '0';
  signal arr1645 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr1645_value\ : value(0 to 67);
  signal \$arr1645_ptr\ : natural range 0 to 99;
  signal \$arr1645_ptr_write\ : natural range 0 to 99;
  signal \$arr1645_write\ : value(0 to 67);
  signal \$arr1645_write_request\ : std_logic := '0';
  signal arr1646 : array_value_72(0 to 99) := (others => (others => '0'));
  signal \$arr1646_value\ : value(0 to 71);
  signal \$arr1646_ptr\ : natural range 0 to 99;
  signal \$arr1646_ptr_write\ : natural range 0 to 99;
  signal \$arr1646_write\ : value(0 to 71);
  signal \$arr1646_write_request\ : std_logic := '0';
  signal arr1647 : array_value_128(0 to 99) := (others => (others => '0'));
  signal \$arr1647_value\ : value(0 to 127);
  signal \$arr1647_ptr\ : natural range 0 to 99;
  signal \$arr1647_ptr_write\ : natural range 0 to 99;
  signal \$arr1647_write\ : value(0 to 127);
  signal \$arr1647_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1643_write_request\ = '1' then
                    arr1643(\$arr1643_ptr_write\) <= \$arr1643_write\;
                  else
                   \$arr1643_value\ <= arr1643(\$arr1643_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1644_write_request\ = '1' then
                    arr1644(\$arr1644_ptr_write\) <= \$arr1644_write\;
                  else
                   \$arr1644_value\ <= arr1644(\$arr1644_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1645_write_request\ = '1' then
                    arr1645(\$arr1645_ptr_write\) <= \$arr1645_write\;
                  else
                   \$arr1645_value\ <= arr1645(\$arr1645_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1646_write_request\ = '1' then
                    arr1646(\$arr1646_ptr_write\) <= \$arr1646_write\;
                  else
                   \$arr1646_value\ <= arr1646(\$arr1646_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr1647_write_request\ = '1' then
                    arr1647(\$arr1647_ptr_write\) <= \$arr1647_write\;
                  else
                   \$arr1647_value\ <= arr1647(\$arr1647_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$136\, \$397\ : value(0 to 1) := (others => '0');
      variable \$144_pow542_arg\, \$146_mul544_arg\, \$147_sub545_arg\, 
               \$402_div543_arg\, \$132_add546_arg\, \$131_sub545_arg\, 
               \$401_pow542_arg\, \$403_mul544_arg\, \$405_add546_arg\, 
               \$128_pow542_arg\, \$129_div543_arg\, \$404_sub545_arg\, 
               \$143_copy_args_to_heap518_arg\, \$145_div543_arg\, 
               \$400_copy_args_to_heap518_arg\, \$148_add546_arg\, 
               \$130_mul544_arg\, \$127_copy_args_to_heap518_arg\ : value(0 to 95) := (others => '0');
      variable \$v1836\, \$v1743\, \$v1818\, \$v1769\, \$v1939\, \$v2077\, 
               \$v2141\, \$v1879\, \$v1717\, \$v2050\, \$v1662\, \$v1829\, 
               \$v1725\, \$v1928\, \$v2133\, \$v1709\, \$v1762\, \$v1890\, 
               \$v1796\, \$v1114\, \$v1766\, \$v2020\, \$v1678\, \$v2027\, 
               \$v1733\, \$v1917\, \$v2003\, \$v1855\, \$v1867\, \$v1807\, 
               \$v1962\, \$v1670\, \$v2149\, \$v1848\, \$v1984\, \$v1901\, 
               \$v1783\, \$v1973\, \$v1950\, \$v2125\, \$v1763\, \$v1686\ : value(0 to 63) := (others => '0');
      variable \$v2093\, \$191_instr\ : value(0 to 71) := (others => '0');
      variable \$v1986\, \$v1809\, \$v1919\, \$v1964\, \$v2052\, \$v1798\, 
               \$v1892\, \$v1975\, \$v1785\, \$v1941\, \$v1881\, \$v1903\, 
               \$v1930\, \$v2216\, \$v1995\, \$v2079\, \$113_p\, p, \$v1820\ : value(0 to 4) := (others => '0');
      variable \$v1996\, \$v1672\, \$v1998\, \$v1802\, \$v2080\, \$v1942\, 
               \$v1664\, \$v1771\, \$v1987\, \$v1789\, \$v2135\, \$v1923\, 
               \$v2053\, \$v1799\, \$v2143\, \$v1896\, \$v1934\, \$v1976\, 
               \$v2022\, \$v1711\, \$v1857\, \$v2083\, \$v1931\, \$v2127\, 
               \$v1885\, \$v1907\, \$v1965\, \$v1920\, \$v1810\, \$v1882\, 
               \$v1850\, \$v1990\, \$v1831\, \$v2094\, \$v1773\, \$v1968\, 
               \$v1735\, \$v1952\, \$v1765\, \$v1945\, \$v1688\, \$v1904\, 
               \$v1680\, \$v2151\, \$v1727\, \$v2056\, \$v1824\, \$v1869\, 
               \$v1719\, \$v1768\, \$v1786\, \$v1893\, \$v1838\, \$v1821\, 
               \$v1979\, \$v1813\, \$v2029\ : value(0 to 3) := (others => '0');
      variable \$149_vm_run_code521_arg\ : value(0 to 294) := (others => '0');
      variable \$v1499\ : value(0 to 127) := (others => '0');
      variable \$v1961\, \$v1685\, \$v1916\, cond, \$v2037\, \$v2139\, 
               \$v2140\, \$v1784\, \$v1938\, \$v1724\, \$v2121\, \$v2107\, 
               \$v2246\, \$v2209\, \$v1828\, rdy1649, condition, \$v1918\, 
               \$v1731\, \$v2123\, \$v1963\, \$v1842\, \$v2231\, \$v2147\, 
               rdy2109, \$v1706\, \$v1747\, \$v1808\, \$v2072\, \$v2199\, 
               \$v2011\, \$v2100\, \$v1988\, \$v2188\, \$v1669\, \$v1940\, x, 
               \$v2098\, \$v1723\, result2108, \$v1693\, \$v1929\, \$v2155\, 
               \$v1862\, \$v1757\, \$v2054\, \$v1668\, \$v1705\, \$v1716\, 
               result2111, \$v1911\, \$v1854\, \$v1684\, \$v2002\, \$v1732\, 
               \$v1782\, \$v1658\, \$v1790\, result1695, \$v1835\, \$v2157\, 
               \$v1878\, \$v2049\, \$v1883\, \$v2099\, \$98_a1\, \$v2051\, 
               \$v1677\, \$v1905\, \$v1707\, \$v2161\, \$v2194\, \$395\, res, 
               \$v1781\, \$v1654\, \$v2204\, \$v2026\, 
               \$149_vm_run_code521_result\, \$v2236\, \$v1739\, \$v2221\, 
               \$v2078\, \$v2102\, \$v1777\, \$v2171\, \$v1866\, \$v1761\, 
               \$v1791\, rdy2112, \$v1787\, result1648, \$v1900\, \$v1660\, 
               \$v1751\, \$v1972\, \$v2132\, \$v1811\, \$v2087\, \$v1974\, 
               \$v1921\, \$v2117\, \$v2081\, rdy1696, \$v2166\, \$v2045\, 
               \$v1932\, \$v2193\, b2, \$v2183\, \$v2041\, \$v2068\, 
               \$v2148\, \$v2033\, \$v2243\, \$v2198\, \$v1822\, \$v1676\, 
               \$115_b\, \$v2244\, \$v1957\, \$v2124\, \$v1708\, \$v1956\, 
               \$v1891\, \$v1795\, \$v1861\, \$v1756\, \$v2177\, \$v1701\, 
               \$v1966\, \$v1902\, \$134_is_loaded\, \$v2092\, \$v1694\, 
               \$v1985\, \$v1741\, \$v2214\, \$v1819\, \$v1994\, \$v1983\, 
               \$v1692\, \$v2060\, \$v2076\, \$v2122\, \$v2226\, \$v1977\, 
               \$v2015\, \$v2088\, \$v1715\, \$v1880\, \$v2131\, \$v1740\, 
               \$v2215\, \$v1817\, \$v2007\, \$v2205\, \$v1797\, \$v1847\, 
               \$v1949\, \$v2019\, \$v1943\, \$v1927\, \$v1800\, \$v2241\, 
               rdy2104, \$v1661\, \$v2237\, \$v1843\, \$v1659\, \$v2156\, 
               \$v1889\, \$v1806\, \$v1894\, \$v1874\, \$v2064\, \$v1873\ : value(0 to 0) := (others => '0');
      variable \$v2210\, \$147_sub545_result\, \$v2222\, fst_operand, 
               \$v2227\, \$511_int_value\, \$631_int_value\, result2103, 
               scd_operand, \$335_divisor\, \$200_i\, base, debut, \$v2189\, 
               \$458_a\, \$482_int_value\, \$99_a\, 
               \$143_copy_args_to_heap518_result\, \$148_add546_result\, 
               \$636_a\, \$v2162\, \$487_a\, \$v2167\, \$353_a\, \$135_cy\, 
               \$114_n\, \$v2172\, \$254_a\, \$196_l\, \$201_i\, 
               \$146_mul544_result\, \$v2184\, \$192_n\, \$283_a\, \$694_a\, 
               \$557_a\, \$195_l\, \$539_divisor\, \$v1752\, \$v1912\, 
               \$307_int_value\, \$193_l\, exponent, \$453_int_value\, 
               \$516_a\, \$v2178\, \$606_int_value\, resultat, 
               \$680_divisor\, \$144_pow542_result\, \$197_i\, 
               \$145_div543_result\, \$312_a\, \$v2232\, \$656_int_value\, 
               \$198_l\, \$199_i\, \$249_int_value\, b, \$278_int_value\, 
               \$393\, \$661_a\, a, \$611_a\ : value(0 to 31) := (others => '0');
      variable \$165\ : value(0 to 293) := (others => '0');
      variable \$v50\, \$v1764\, \$v124\, \$v1944\, \$v1726\, \$v1989\, 
               \$v142\, \$v229\, \$v2217\, \$v1837\, \$v159\, \$v149\, 
               \$v1884\, \$v2028\, \$v1997\, second_value, \$v56\, \$452_v\, 
               first_value, \$352\, \$v187\, \$v221\, \$248_v\, \$v184\, 
               \$v1823\, \$v2142\, \$v2055\, \$v1951\, \$389\, \$655_v\, 
               \$v1967\, \$v1767\, \$v47\, \$v66\, \$v1663\, \$v45\, 
               \$v1978\, \$306_v\, \$v92\, \$v225\, \$630_v\, var, \$v2150\, 
               \$v68\, \$v1742\, \$v1906\, \$v1679\, \$v1770\, \$726\, 
               \$v1801\, \$v114\, \$693\, \$v1812\, \$v1856\, \$v1830\, 
               \$v1933\, \$556\, \$v194\, \$v1772\, \$v1687\, \$v1895\, 
               \value\, \$v2126\, \$v2179\, \$v1868\, \$v1710\, \$v1788\, 
               \$v152\, \$v237\, \$v2082\, \$v1671\, \$v117\, \$v1849\, 
               \$277_v\, \$481_v\, \$v2173\, \$v2200\, \$204_v\, \$593\, 
               \$v1718\, local_value, \$v2021\, \$v1922\, \$v2134\, \$v1734\, 
               \$v53\, v, \$510_v\, \$605_v\ : value(0 to 67) := (others => '0');
      variable \$arr1643_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1644_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1645_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1646_ptr_take\ : value(0 to 0) := "0";
      variable \$arr1647_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(\$611_a\); default_zero(\$v1873\); default_zero(a); 
          default_zero(\$v1686\); default_zero(\$605_v\); 
          default_zero(\$v2064\); default_zero(\$661_a\); 
          default_zero(\$v2029\); default_zero(\$v1874\); 
          default_zero(\$v1894\); 
          default_zero(\$127_copy_args_to_heap518_arg\); 
          default_zero(\$v1763\); default_zero(\$v1806\); 
          default_zero(\$393\); default_zero(\$v2125\); 
          default_zero(\$v1889\); default_zero(\$v1813\); 
          default_zero(\$v2156\); default_zero(\$v1659\); 
          default_zero(\$v1843\); default_zero(\$510_v\); 
          default_zero(\$v2237\); default_zero(\$v1661\); default_zero(v); 
          default_zero(rdy2104); default_zero(\$v2241\); 
          default_zero(\$v1950\); default_zero(\$278_int_value\); 
          default_zero(\$v53\); default_zero(\$130_mul544_arg\); 
          default_zero(\$v1800\); default_zero(\$v1734\); 
          default_zero(\$v1973\); default_zero(\$397\); 
          default_zero(\$v1927\); default_zero(\$v1783\); 
          default_zero(\$v1943\); default_zero(b); 
          default_zero(\$148_add546_arg\); default_zero(\$v1979\); 
          default_zero(\$v2019\); default_zero(\$v1901\); 
          default_zero(\$249_int_value\); default_zero(\$v2134\); 
          default_zero(\$v1949\); default_zero(\$v1847\); 
          default_zero(\$v1797\); default_zero(\$v1922\); 
          default_zero(\$400_copy_args_to_heap518_arg\); 
          default_zero(\$199_i\); default_zero(\$v2021\); 
          default_zero(\$v2205\); default_zero(\$v1984\); 
          default_zero(local_value); default_zero(\$v1821\); 
          default_zero(\$198_l\); default_zero(\$v1718\); 
          default_zero(\$145_div543_arg\); default_zero(\$v2007\); 
          default_zero(\$593\); default_zero(\$v1838\); 
          default_zero(\$v1817\); default_zero(\$656_int_value\); 
          default_zero(\$v2215\); default_zero(\$v1893\); 
          default_zero(\$v1740\); default_zero(\$v1848\); 
          default_zero(\$v2131\); default_zero(\$v1880\); 
          default_zero(\$204_v\); default_zero(\$v2232\); 
          default_zero(\$143_copy_args_to_heap518_arg\); 
          default_zero(\$v2200\); default_zero(\$312_a\); 
          default_zero(\$145_div543_result\); default_zero(\$197_i\); 
          default_zero(\$v2173\); default_zero(\$481_v\); 
          default_zero(\$v1715\); default_zero(\$277_v\); 
          default_zero(\$v2088\); default_zero(\$v2015\); 
          default_zero(\$v1977\); default_zero(\$v2226\); 
          default_zero(\$v2122\); default_zero(\$v2076\); 
          default_zero(\$v2060\); default_zero(\$v1849\); 
          default_zero(\$144_pow542_result\); default_zero(\$v1692\); 
          default_zero(\$v2149\); default_zero(\$v117\); 
          default_zero(\$v1670\); default_zero(\$v1786\); 
          default_zero(\$v1983\); default_zero(\$v1768\); 
          default_zero(\$v1994\); default_zero(\$v1819\); 
          default_zero(\$680_divisor\); default_zero(resultat); 
          default_zero(\$149_vm_run_code521_arg\); 
          default_zero(\$606_int_value\); default_zero(\$v2214\); 
          default_zero(\$v1719\); default_zero(\$v1869\); 
          default_zero(\$v1499\); default_zero(\$v1824\); 
          default_zero(\$v1671\); default_zero(\$v1741\); 
          default_zero(\$v1985\); default_zero(\$v2082\); 
          default_zero(\$v1694\); default_zero(\$v1962\); 
          default_zero(\$v2178\); default_zero(\$516_a\); 
          default_zero(\$v2092\); default_zero(\$134_is_loaded\); 
          default_zero(\$v1902\); default_zero(\$v237\); 
          default_zero(\$v1807\); default_zero(\$v1966\); 
          default_zero(\$v152\); default_zero(\$v1701\); 
          default_zero(\$v2177\); default_zero(\$453_int_value\); 
          default_zero(\$v1756\); default_zero(\$v2056\); 
          default_zero(\$v1867\); default_zero(\$v1788\); 
          default_zero(\$v1861\); default_zero(\$v1727\); 
          default_zero(\$404_sub545_arg\); default_zero(\$v1795\); 
          default_zero(\$v1820\); default_zero(exponent); 
          default_zero(\$v1891\); default_zero(\$v1710\); 
          default_zero(\$129_div543_arg\); default_zero(\$v1868\); 
          default_zero(\$v2179\); default_zero(\$v2126\); 
          default_zero(\$193_l\); default_zero(p); default_zero(\$v1956\); 
          default_zero(\value\); default_zero(\$v1855\); 
          default_zero(\$v2151\); default_zero(\$v1708\); 
          default_zero(\$v1680\); default_zero(\$v2124\); 
          default_zero(\$v1957\); default_zero(\$v1895\); 
          default_zero(\$v2244\); default_zero(\$115_b\); 
          default_zero(\$v1687\); default_zero(\$307_int_value\); 
          default_zero(\$v1676\); default_zero(\$v1772\); 
          default_zero(\$v1904\); default_zero(\$v1822\); 
          default_zero(\$v2198\); default_zero(\$v2243\); 
          default_zero(\$v1688\); default_zero(\$v2033\); 
          default_zero(\$v2148\); default_zero(\$v2003\); 
          default_zero(\$113_p\); default_zero(\$v1912\); 
          default_zero(\$v2068\); default_zero(\$v194\); 
          default_zero(\$v1752\); default_zero(\$556\); 
          default_zero(\$v1933\); default_zero(\$v1945\); 
          default_zero(\$v1765\); default_zero(\$v2041\); 
          default_zero(\$v1830\); default_zero(\$v2183\); 
          default_zero(\$v1856\); default_zero(\$v1812\); 
          default_zero(\$693\); default_zero(\$128_pow542_arg\); 
          default_zero(\$v114\); default_zero(\$539_divisor\); 
          default_zero(\$v1952\); default_zero(b2); default_zero(\$v2193\); 
          default_zero(\$195_l\); default_zero(\$v1932\); 
          default_zero(\$v1801\); default_zero(\$v2045\); 
          default_zero(\$v2166\); default_zero(rdy1696); 
          default_zero(\$557_a\); default_zero(\$v1917\); 
          default_zero(\$v1735\); default_zero(\$694_a\); 
          default_zero(\$v2081\); default_zero(\$v2117\); 
          default_zero(\$v1921\); default_zero(\$405_add546_arg\); 
          default_zero(\$726\); default_zero(\$v1974\); 
          default_zero(\$283_a\); default_zero(\$v2087\); 
          default_zero(\$v1811\); default_zero(\$v2132\); 
          default_zero(\$v1972\); default_zero(\$v1770\); 
          default_zero(\$v1733\); default_zero(\$v1751\); 
          default_zero(\$v1679\); default_zero(\$v2027\); 
          default_zero(\$v1968\); default_zero(\$v1660\); 
          default_zero(\$192_n\); default_zero(\$v1900\); 
          default_zero(\$v1906\); default_zero(\$v1742\); 
          default_zero(result1648); default_zero(\$v1787\); 
          default_zero(rdy2112); default_zero(\$v1791\); 
          default_zero(\$v1678\); default_zero(\$v1761\); 
          default_zero(\$v1773\); default_zero(\$v2184\); 
          default_zero(\$146_mul544_result\); default_zero(\$v2094\); 
          default_zero(\$201_i\); default_zero(\$v68\); 
          default_zero(\$v1866\); default_zero(\$v2150\); 
          default_zero(\$v2171\); default_zero(\$v1831\); 
          default_zero(\$v1777\); default_zero(var); default_zero(\$630_v\); 
          default_zero(\$v2020\); default_zero(\$v2102\); 
          default_zero(\$v225\); default_zero(\$196_l\); 
          default_zero(\$v2078\); default_zero(\$254_a\); 
          default_zero(\$v2221\); default_zero(\$v1739\); 
          default_zero(\$v1990\); default_zero(\$v1850\); 
          default_zero(\$v2236\); default_zero(\$v2172\); 
          default_zero(\$v1882\); default_zero(\$v1810\); 
          default_zero(\$114_n\); default_zero(\$135_cy\); 
          default_zero(\$353_a\); default_zero(\$191_instr\); 
          default_zero(\$v92\); default_zero(\$149_vm_run_code521_result\); 
          default_zero(\$v1920\); default_zero(\$v2026\); 
          default_zero(\$v1965\); default_zero(\$v1907\); 
          default_zero(\$v2167\); default_zero(\$v1885\); 
          default_zero(\$306_v\); default_zero(\$v2204\); 
          default_zero(\$487_a\); default_zero(\$v2127\); 
          default_zero(\$v1654\); default_zero(\$v2079\); 
          default_zero(\$v1781\); default_zero(\$v1978\); default_zero(res); 
          default_zero(\$395\); default_zero(\$v2194\); 
          default_zero(\$v2161\); default_zero(\$v1707\); 
          default_zero(\$v1905\); default_zero(\$v1766\); 
          default_zero(\$v1931\); default_zero(\$v1677\); 
          default_zero(\$v2083\); default_zero(\$v1995\); 
          default_zero(\$403_mul544_arg\); default_zero(\$v1114\); 
          default_zero(\$v2051\); default_zero(\$v1857\); 
          default_zero(\$98_a1\); default_zero(\$v2162\); 
          default_zero(\$636_a\); default_zero(\$v45\); 
          default_zero(\$v2099\); default_zero(\$v1711\); 
          default_zero(\$v1883\); default_zero(\$v2216\); 
          default_zero(\$v2022\); default_zero(\$148_add546_result\); 
          default_zero(\$v1930\); default_zero(\$v2049\); 
          default_zero(\$v1878\); 
          default_zero(\$143_copy_args_to_heap518_result\); 
          default_zero(\$v1663\); default_zero(\$v2157\); 
          default_zero(\$v1835\); default_zero(result1695); 
          default_zero(\$v1790\); default_zero(\$v66\); 
          default_zero(\$v1658\); default_zero(\$v1796\); 
          default_zero(\$v1782\); default_zero(\$v47\); 
          default_zero(\$v1890\); default_zero(\$v1767\); 
          default_zero(\$v1732\); default_zero(\$v1967\); 
          default_zero(\$v1762\); default_zero(\$v2002\); 
          default_zero(\$v1709\); default_zero(\$v2133\); 
          default_zero(\$v1976\); default_zero(\$655_v\); 
          default_zero(\$v1684\); default_zero(\$389\); 
          default_zero(\$v1934\); default_zero(\$v1854\); 
          default_zero(\$99_a\); default_zero(\$v1911\); 
          default_zero(result2111); default_zero(\$v1928\); 
          default_zero(\$v1716\); default_zero(\$v1951\); 
          default_zero(\$v1705\); default_zero(\$v1668\); 
          default_zero(\$v1725\); default_zero(\$v2054\); 
          default_zero(\$v1757\); default_zero(\$v1896\); 
          default_zero(\$v1829\); default_zero(\$482_int_value\); 
          default_zero(\$v1862\); default_zero(\$v2155\); 
          default_zero(\$v2143\); default_zero(\$v1929\); 
          default_zero(\$v1693\); default_zero(result2108); 
          default_zero(\$v2055\); default_zero(\$v1723\); 
          default_zero(\$v2142\); default_zero(\$v1662\); 
          default_zero(\$v2098\); default_zero(\$401_pow542_arg\); 
          default_zero(x); default_zero(\$v1799\); default_zero(\$v1940\); 
          default_zero(\$v1823\); default_zero(\$v1669\); 
          default_zero(\$v184\); default_zero(\$v2188\); 
          default_zero(\$v1988\); default_zero(\$248_v\); 
          default_zero(\$458_a\); default_zero(\$136\); 
          default_zero(\$v2189\); default_zero(\$131_sub545_arg\); 
          default_zero(\$v2053\); default_zero(\$v1903\); 
          default_zero(\$v221\); default_zero(debut); 
          default_zero(\$132_add546_arg\); default_zero(\$v187\); 
          default_zero(\$v1881\); default_zero(\$v1923\); 
          default_zero(\$v1941\); default_zero(\$v2100\); 
          default_zero(\$v2011\); default_zero(\$352\); default_zero(\$165\); 
          default_zero(\$v2199\); default_zero(base); default_zero(\$v2135\); 
          default_zero(\$v1789\); default_zero(first_value); 
          default_zero(\$v2050\); default_zero(\$v1785\); 
          default_zero(\$200_i\); default_zero(\$v2072\); 
          default_zero(\$v1808\); default_zero(\$335_divisor\); 
          default_zero(\$v1747\); default_zero(\$v1987\); 
          default_zero(\$v1706\); default_zero(\$v1717\); 
          default_zero(\$452_v\); default_zero(\$v1975\); 
          default_zero(rdy2109); default_zero(\$v56\); 
          default_zero(\$v1892\); default_zero(scd_operand); 
          default_zero(second_value); default_zero(\$v2147\); 
          default_zero(\$v2231\); default_zero(\$v1771\); 
          default_zero(\$402_div543_arg\); default_zero(\$v1997\); 
          default_zero(\$v2028\); default_zero(result2103); 
          default_zero(\$v1879\); default_zero(\$631_int_value\); 
          default_zero(\$v1842\); default_zero(\$v1664\); 
          default_zero(\$v1942\); default_zero(\$511_int_value\); 
          default_zero(\$v1884\); default_zero(\$v1798\); 
          default_zero(\$v1963\); default_zero(\$147_sub545_arg\); 
          default_zero(\$v2123\); default_zero(\$146_mul544_arg\); 
          default_zero(\$v2141\); default_zero(\$v149\); 
          default_zero(\$v1731\); default_zero(\$v159\); 
          default_zero(\$v2227\); default_zero(\$v1837\); 
          default_zero(\$v2080\); default_zero(\$v1918\); 
          default_zero(condition); default_zero(fst_operand); 
          default_zero(\$v2052\); default_zero(\$v2217\); 
          default_zero(\$v229\); default_zero(\$v1802\); 
          default_zero(rdy1649); default_zero(\$v2093\); 
          default_zero(\$v2077\); default_zero(\$v2222\); 
          default_zero(\$v142\); default_zero(\$v1828\); 
          default_zero(\$v2209\); default_zero(\$v1989\); 
          default_zero(\$v2246\); default_zero(\$v2107\); 
          default_zero(\$v1939\); default_zero(\$v2121\); 
          default_zero(\$147_sub545_result\); default_zero(\$v1769\); 
          default_zero(\$v1998\); default_zero(\$v1964\); 
          default_zero(\$v1726\); default_zero(\$v1724\); 
          default_zero(\$v1672\); default_zero(\$v1944\); 
          default_zero(\$v2210\); default_zero(\$v1938\); 
          default_zero(\$v1919\); default_zero(\$v1818\); 
          default_zero(\$v1743\); default_zero(\$v1784\); 
          default_zero(\$v2140\); default_zero(\$v1809\); 
          default_zero(\$v1986\); default_zero(\$v124\); 
          default_zero(\$v2139\); default_zero(\$v2037\); default_zero(cond); 
          default_zero(\$v1836\); default_zero(\$v1764\); 
          default_zero(\$v1916\); default_zero(\$v1685\); 
          default_zero(\$v50\); default_zero(\$v1996\); 
          default_zero(\$v1961\); default_zero(\$144_pow542_arg\); 
          rdy <= "1";
          rdy1649 := "0";
          \state\ <= compute1650;
          state_var2250 <= compute2113;
          state_var2249 <= compute2110;
          state_var2248 <= compute2105;
          state_var2247 <= compute1697;
          
        else if run = '1' then
          case \state\ is
          when \$127_copy_args_to_heap518\ =>
            \$v1659\ := eclat_eq(\$127_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1659\(0) = '1' then
              \state\ <= \$127_copy_args_to_heap518\;
            else
              \$v1658\ := \$arr1644_ptr_take\;
              if \$v1658\(0) = '1' then
                \state\ <= q_wait1657;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$127_copy_args_to_heap518_arg\(32 to 63) & \$127_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
                \state\ <= pause_getI1655;
              end if;
            end if;
          when \$128_pow542\ =>
            \$v1660\ := eclat_eq(\$128_pow542_arg\(32 to 63) & "00000000000000000000000000000000");
            if \$v1660\(0) = '1' then
              \state\ <= \$128_pow542\;
            else
              \$128_pow542_arg\ := \$128_pow542_arg\(0 to 31) & eclat_sub(\$128_pow542_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$128_pow542_arg\(64 to 95) & \$128_pow542_arg\(0 to 31));
              \state\ <= \$128_pow542\;
            end if;
          when \$129_div543\ =>
            \$v1669\ := eclat_eq(\$129_div543_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1669\(0) = '1' then
              \state\ <= \$129_div543\;
            else
              \$v1668\ := \$arr1644_ptr_take\;
              if \$v1668\(0) = '1' then
                \state\ <= q_wait1667;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$129_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$129_div543_arg\(0 to 31))));
                \state\ <= pause_getI1665;
              end if;
            end if;
          when \$130_mul544\ =>
            \$v1677\ := eclat_eq(\$130_mul544_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1677\(0) = '1' then
              \state\ <= \$130_mul544\;
            else
              \$v1676\ := \$arr1644_ptr_take\;
              if \$v1676\(0) = '1' then
                \state\ <= q_wait1675;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_mul544_arg\(0 to 31))));
                \state\ <= pause_getI1673;
              end if;
            end if;
          when \$131_sub545\ =>
            \$v1685\ := eclat_eq(\$131_sub545_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1685\(0) = '1' then
              \state\ <= \$131_sub545\;
            else
              \$v1684\ := \$arr1644_ptr_take\;
              if \$v1684\(0) = '1' then
                \state\ <= q_wait1683;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_sub545_arg\(0 to 31))));
                \state\ <= pause_getI1681;
              end if;
            end if;
          when \$132_add546\ =>
            \$v1693\ := eclat_eq(\$132_add546_arg\(0 to 31) & "00000000000000000000000000000000");
            if \$v1693\(0) = '1' then
              \state\ <= \$132_add546\;
            else
              \$v1692\ := \$arr1644_ptr_take\;
              if \$v1692\(0) = '1' then
                \state\ <= q_wait1691;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_add546_arg\(0 to 31))));
                \state\ <= pause_getI1689;
              end if;
            end if;
          when \$615_forever5481612\ =>
            \state\ <= \$615_forever5481612\;
          when \$640_forever5481611\ =>
            \state\ <= \$640_forever5481611\;
          when \$665_forever5481610\ =>
            \state\ <= \$665_forever5481610\;
          when \$689_forever5481608\ =>
            \state\ <= \$689_forever5481608\;
          when \$698_forever5481609\ =>
            \state\ <= \$698_forever5481609\;
          when pause_getI1655 =>
            \state\ <= pause_getII1656;
          when pause_getI1665 =>
            \state\ <= pause_getII1666;
          when pause_getI1673 =>
            \state\ <= pause_getII1674;
          when pause_getI1681 =>
            \state\ <= pause_getII1682;
          when pause_getI1689 =>
            \state\ <= pause_getII1690;
          when pause_getII1656 =>
            \$arr1644_ptr_take\(0) := '0';
            \$726\ := \$arr1644_value\;
            \$v1654\ := \$arr1643_ptr_take\;
            if \$v1654\(0) = '1' then
              \state\ <= q_wait1653;
            else
              \$arr1643_ptr_take\(0) := '1';
              \$arr1643_ptr_write\ <= to_integer(unsigned(\$127_copy_args_to_heap518_arg\(64 to 95)));
              \$arr1643_write_request\ <= '1';
              \$arr1643_write\ <= \$726\;
              \state\ <= pause_setI1651;
            end if;
          when pause_getII1666 =>
            \$arr1644_ptr_take\(0) := '0';
            \$693\ := \$arr1644_value\;
            \$v1663\ := \$693\;
            \$v1664\ := \$v1663\(0 to 3);
            \$v1662\ := \$v1663\(4 to 67);
            case \$v1664\ is
            when "0001" =>
              \$694_a\ := \$v1662\(0 to 31);
              \$680_divisor\ := \$694_a\;
              \$v1661\ := eclat_eq(\$680_divisor\ & "00000000000000000000000000000000");
              if \$v1661\(0) = '1' then
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("Division par zero"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$689_forever5481608\;
              else
                \$129_div543_arg\ := eclat_sub(\$129_div543_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$129_div543_arg\(32 to 63) & \$680_divisor\) & \$129_div543_arg\(64 to 95);
                \state\ <= \$129_div543\;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$698_forever5481609\;
            end case;
          when pause_getII1674 =>
            \$arr1644_ptr_take\(0) := '0';
            \$655_v\ := \$arr1644_value\;
            \$v1671\ := \$655_v\;
            \$v1672\ := \$v1671\(0 to 3);
            \$v1670\ := \$v1671\(4 to 67);
            case \$v1672\ is
            when "0001" =>
              \$661_a\ := \$v1670\(0 to 31);
              \$656_int_value\ := \$661_a\;
              \$130_mul544_arg\ := eclat_sub(\$130_mul544_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$130_mul544_arg\(32 to 63) & \$656_int_value\) & \$130_mul544_arg\(64 to 95);
              \state\ <= \$130_mul544\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$665_forever5481610\;
            end case;
          when pause_getII1682 =>
            \$arr1644_ptr_take\(0) := '0';
            \$630_v\ := \$arr1644_value\;
            \$v1679\ := \$630_v\;
            \$v1680\ := \$v1679\(0 to 3);
            \$v1678\ := \$v1679\(4 to 67);
            case \$v1680\ is
            when "0001" =>
              \$636_a\ := \$v1678\(0 to 31);
              \$631_int_value\ := \$636_a\;
              \$131_sub545_arg\ := eclat_sub(\$131_sub545_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$131_sub545_arg\(32 to 63) & \$631_int_value\) & \$131_sub545_arg\(64 to 95);
              \state\ <= \$131_sub545\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$640_forever5481611\;
            end case;
          when pause_getII1690 =>
            \$arr1644_ptr_take\(0) := '0';
            \$605_v\ := \$arr1644_value\;
            \$v1687\ := \$605_v\;
            \$v1688\ := \$v1687\(0 to 3);
            \$v1686\ := \$v1687\(4 to 67);
            case \$v1688\ is
            when "0001" =>
              \$611_a\ := \$v1686\(0 to 31);
              \$606_int_value\ := \$611_a\;
              \$132_add546_arg\ := eclat_sub(\$132_add546_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$132_add546_arg\(32 to 63) & \$606_int_value\) & \$132_add546_arg\(64 to 95);
              \state\ <= \$132_add546\;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$615_forever5481612\;
            end case;
          when pause_setI1651 =>
            \$arr1643_write_request\ <= '0';
            \state\ <= pause_setII1652;
          when pause_setII1652 =>
            \$arr1643_ptr_take\(0) := '0';
            \$127_copy_args_to_heap518_arg\ := eclat_sub(\$127_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000001") & \$127_copy_args_to_heap518_arg\(32 to 63) & eclat_add(\$127_copy_args_to_heap518_arg\(64 to 95) & "00000000000000000000000000000001");
            \state\ <= \$127_copy_args_to_heap518\;
          when q_wait1653 =>
            \$v1654\ := \$arr1643_ptr_take\;
            if \$v1654\(0) = '1' then
              \state\ <= q_wait1653;
            else
              \$arr1643_ptr_take\(0) := '1';
              \$arr1643_ptr_write\ <= to_integer(unsigned(\$127_copy_args_to_heap518_arg\(64 to 95)));
              \$arr1643_write_request\ <= '1';
              \$arr1643_write\ <= \$726\;
              \state\ <= pause_setI1651;
            end if;
          when q_wait1657 =>
            \$v1658\ := \$arr1644_ptr_take\;
            if \$v1658\(0) = '1' then
              \state\ <= q_wait1657;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$127_copy_args_to_heap518_arg\(32 to 63) & \$127_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI1655;
            end if;
          when q_wait1667 =>
            \$v1668\ := \$arr1644_ptr_take\;
            if \$v1668\(0) = '1' then
              \state\ <= q_wait1667;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$129_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$129_div543_arg\(0 to 31))));
              \state\ <= pause_getI1665;
            end if;
          when q_wait1675 =>
            \$v1676\ := \$arr1644_ptr_take\;
            if \$v1676\(0) = '1' then
              \state\ <= q_wait1675;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$130_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$130_mul544_arg\(0 to 31))));
              \state\ <= pause_getI1673;
            end if;
          when q_wait1683 =>
            \$v1684\ := \$arr1644_ptr_take\;
            if \$v1684\(0) = '1' then
              \state\ <= q_wait1683;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$131_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$131_sub545_arg\(0 to 31))));
              \state\ <= pause_getI1681;
            end if;
          when q_wait1691 =>
            \$v1692\ := \$arr1644_ptr_take\;
            if \$v1692\(0) = '1' then
              \state\ <= q_wait1691;
            else
              \$arr1644_ptr_take\(0) := '1';
              \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$132_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$132_add546_arg\(0 to 31))));
              \state\ <= pause_getI1689;
            end if;
          when compute1650 =>
            rdy1649 := eclat_false;
            case state_var2249 is
            when compute2110 =>
              rdy2109 := eclat_false;
              \$v2244\ := \$395\;
              if \$v2244\(0) = '1' then
                result2108 := eclat_true;
                rdy2109 := eclat_true;
                state_var2249 <= compute2110;
              else
                case state_var2250 is
                when \$400_copy_args_to_heap518\ =>
                  \$v2122\ := eclat_eq(\$400_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2122\(0) = '1' then
                    state_var2250 <= \$400_copy_args_to_heap518\;
                  else
                    \$v2121\ := \$arr1644_ptr_take\;
                    if \$v2121\(0) = '1' then
                      state_var2250 <= q_wait2120;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$400_copy_args_to_heap518_arg\(32 to 63) & \$400_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
                      state_var2250 <= pause_getI2118;
                    end if;
                  end if;
                when \$401_pow542\ =>
                  \$v2123\ := eclat_eq(\$401_pow542_arg\(32 to 63) & "00000000000000000000000000000000");
                  if \$v2123\(0) = '1' then
                    state_var2250 <= \$401_pow542\;
                  else
                    \$401_pow542_arg\ := \$401_pow542_arg\(0 to 31) & eclat_sub(\$401_pow542_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$401_pow542_arg\(64 to 95) & \$401_pow542_arg\(0 to 31));
                    state_var2250 <= \$401_pow542\;
                  end if;
                when \$402_div543\ =>
                  \$v2132\ := eclat_eq(\$402_div543_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2132\(0) = '1' then
                    state_var2250 <= \$402_div543\;
                  else
                    \$v2131\ := \$arr1644_ptr_take\;
                    if \$v2131\(0) = '1' then
                      state_var2250 <= q_wait2130;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$402_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$402_div543_arg\(0 to 31))));
                      state_var2250 <= pause_getI2128;
                    end if;
                  end if;
                when \$403_mul544\ =>
                  \$v2140\ := eclat_eq(\$403_mul544_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2140\(0) = '1' then
                    state_var2250 <= \$403_mul544\;
                  else
                    \$v2139\ := \$arr1644_ptr_take\;
                    if \$v2139\(0) = '1' then
                      state_var2250 <= q_wait2138;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$403_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$403_mul544_arg\(0 to 31))));
                      state_var2250 <= pause_getI2136;
                    end if;
                  end if;
                when \$404_sub545\ =>
                  \$v2148\ := eclat_eq(\$404_sub545_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2148\(0) = '1' then
                    state_var2250 <= \$404_sub545\;
                  else
                    \$v2147\ := \$arr1644_ptr_take\;
                    if \$v2147\(0) = '1' then
                      state_var2250 <= q_wait2146;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$404_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$404_sub545_arg\(0 to 31))));
                      state_var2250 <= pause_getI2144;
                    end if;
                  end if;
                when \$405_add546\ =>
                  \$v2156\ := eclat_eq(\$405_add546_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v2156\(0) = '1' then
                    state_var2250 <= \$405_add546\;
                  else
                    \$v2155\ := \$arr1644_ptr_take\;
                    if \$v2155\(0) = '1' then
                      state_var2250 <= q_wait2154;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$405_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$405_add546_arg\(0 to 31))));
                      state_var2250 <= pause_getI2152;
                    end if;
                  end if;
                when \$462_forever5481642\ =>
                  state_var2250 <= \$466_forever5481636\;
                when \$466_forever5481636\ =>
                  state_var2250 <= \$466_forever5481636\;
                when \$491_forever5481641\ =>
                  state_var2250 <= \$495_forever5481636\;
                when \$495_forever5481636\ =>
                  state_var2250 <= \$495_forever5481636\;
                when \$520_forever5481640\ =>
                  state_var2250 <= \$524_forever5481636\;
                when \$524_forever5481636\ =>
                  state_var2250 <= \$524_forever5481636\;
                when \$548_forever5481638\ =>
                  state_var2250 <= \$552_forever5481636\;
                when \$552_forever5481636\ =>
                  state_var2250 <= \$552_forever5481636\;
                when \$561_forever5481639\ =>
                  state_var2250 <= \$565_forever5481636\;
                when \$565_forever5481636\ =>
                  state_var2250 <= \$565_forever5481636\;
                when pause_getI2118 =>
                  state_var2250 <= pause_getII2119;
                when pause_getI2128 =>
                  state_var2250 <= pause_getII2129;
                when pause_getI2136 =>
                  state_var2250 <= pause_getII2137;
                when pause_getI2144 =>
                  state_var2250 <= pause_getII2145;
                when pause_getI2152 =>
                  state_var2250 <= pause_getII2153;
                when pause_getII2119 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$593\ := \$arr1644_value\;
                  \$v2117\ := \$arr1643_ptr_take\;
                  if \$v2117\(0) = '1' then
                    state_var2250 <= q_wait2116;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr_write\ <= to_integer(unsigned(\$400_copy_args_to_heap518_arg\(64 to 95)));
                    \$arr1643_write_request\ <= '1';
                    \$arr1643_write\ <= \$593\;
                    state_var2250 <= pause_setI2114;
                  end if;
                when pause_getII2129 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$556\ := \$arr1644_value\;
                  \$v2126\ := \$556\;
                  \$v2127\ := \$v2126\(0 to 3);
                  \$v2125\ := \$v2126\(4 to 67);
                  case \$v2127\ is
                  when "0001" =>
                    \$557_a\ := \$v2125\(0 to 31);
                    \$539_divisor\ := \$557_a\;
                    \$v2124\ := eclat_eq(\$539_divisor\ & "00000000000000000000000000000000");
                    if \$v2124\(0) = '1' then
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("Division par zero"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var2250 <= \$548_forever5481638\;
                    else
                      \$402_div543_arg\ := eclat_sub(\$402_div543_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$402_div543_arg\(32 to 63) & \$539_divisor\) & \$402_div543_arg\(64 to 95);
                      state_var2250 <= \$402_div543\;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2250 <= \$561_forever5481639\;
                  end case;
                when pause_getII2137 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$510_v\ := \$arr1644_value\;
                  \$v2134\ := \$510_v\;
                  \$v2135\ := \$v2134\(0 to 3);
                  \$v2133\ := \$v2134\(4 to 67);
                  case \$v2135\ is
                  when "0001" =>
                    \$516_a\ := \$v2133\(0 to 31);
                    \$511_int_value\ := \$516_a\;
                    \$403_mul544_arg\ := eclat_sub(\$403_mul544_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$403_mul544_arg\(32 to 63) & \$511_int_value\) & \$403_mul544_arg\(64 to 95);
                    state_var2250 <= \$403_mul544\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2250 <= \$520_forever5481640\;
                  end case;
                when pause_getII2145 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$481_v\ := \$arr1644_value\;
                  \$v2142\ := \$481_v\;
                  \$v2143\ := \$v2142\(0 to 3);
                  \$v2141\ := \$v2142\(4 to 67);
                  case \$v2143\ is
                  when "0001" =>
                    \$487_a\ := \$v2141\(0 to 31);
                    \$482_int_value\ := \$487_a\;
                    \$404_sub545_arg\ := eclat_sub(\$404_sub545_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$404_sub545_arg\(32 to 63) & \$482_int_value\) & \$404_sub545_arg\(64 to 95);
                    state_var2250 <= \$404_sub545\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2250 <= \$491_forever5481641\;
                  end case;
                when pause_getII2153 =>
                  \$arr1644_ptr_take\(0) := '0';
                  \$452_v\ := \$arr1644_value\;
                  \$v2150\ := \$452_v\;
                  \$v2151\ := \$v2150\(0 to 3);
                  \$v2149\ := \$v2150\(4 to 67);
                  case \$v2151\ is
                  when "0001" =>
                    \$458_a\ := \$v2149\(0 to 31);
                    \$453_int_value\ := \$458_a\;
                    \$405_add546_arg\ := eclat_sub(\$405_add546_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$405_add546_arg\(32 to 63) & \$453_int_value\) & \$405_add546_arg\(64 to 95);
                    state_var2250 <= \$405_add546\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2250 <= \$462_forever5481642\;
                  end case;
                when pause_setI2114 =>
                  \$arr1643_write_request\ <= '0';
                  state_var2250 <= pause_setII2115;
                when pause_setI2158 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2159;
                when pause_setI2163 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2164;
                when pause_setI2168 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2169;
                when pause_setI2174 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2175;
                when pause_setI2180 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2181;
                when pause_setI2185 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2186;
                when pause_setI2190 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2191;
                when pause_setI2195 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2196;
                when pause_setI2201 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2202;
                when pause_setI2206 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2207;
                when pause_setI2211 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2212;
                when pause_setI2218 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2219;
                when pause_setI2223 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2224;
                when pause_setI2228 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2229;
                when pause_setI2233 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2234;
                when pause_setI2238 =>
                  \$arr1646_write_request\ <= '0';
                  state_var2250 <= pause_setII2239;
                when pause_setII2115 =>
                  \$arr1643_ptr_take\(0) := '0';
                  \$400_copy_args_to_heap518_arg\ := eclat_sub(\$400_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000001") & \$400_copy_args_to_heap518_arg\(32 to 63) & eclat_add(\$400_copy_args_to_heap518_arg\(64 to 95) & "00000000000000000000000000000001");
                  state_var2250 <= \$400_copy_args_to_heap518\;
                when pause_setII2159 =>
                  \$arr1646_ptr_take\(0) := '0';
                  result2111 := eclat_unit;
                  rdy2112 := eclat_true;
                  state_var2250 <= compute2113;
                when pause_setII2164 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2161\ := \$arr1646_ptr_take\;
                  if \$v2161\(0) = '1' then
                    state_var2250 <= q_wait2160;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2157\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 15;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0111" & \$v2157\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2158;
                  end if;
                when pause_setII2169 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2166\ := \$arr1646_ptr_take\;
                  if \$v2166\(0) = '1' then
                    state_var2250 <= q_wait2165;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2162\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 14;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2162\&X"000000000";
                    state_var2250 <= pause_setI2163;
                  end if;
                when pause_setII2175 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2171\ := \$arr1646_ptr_take\;
                  if \$v2171\(0) = '1' then
                    state_var2250 <= q_wait2170;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2167\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 13;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0010" & \$v2167\&X"000000000";
                    state_var2250 <= pause_setI2168;
                  end if;
                when pause_setII2181 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2177\ := \$arr1646_ptr_take\;
                  if \$v2177\(0) = '1' then
                    state_var2250 <= q_wait2176;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2172\ := "00000000000000000000000000000001";
                    \$v2173\ := "0001" & \$v2172\&X"00000000";
                    \$arr1646_ptr_write\ <= 12;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2173\;
                    state_var2250 <= pause_setI2174;
                  end if;
                when pause_setII2186 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2183\ := \$arr1646_ptr_take\;
                  if \$v2183\(0) = '1' then
                    state_var2250 <= q_wait2182;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2178\ := "00000000000000000000000000000010";
                    \$v2179\ := "0001" & \$v2178\&X"00000000";
                    \$arr1646_ptr_write\ <= 11;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2179\;
                    state_var2250 <= pause_setI2180;
                  end if;
                when pause_setII2191 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2188\ := \$arr1646_ptr_take\;
                  if \$v2188\(0) = '1' then
                    state_var2250 <= q_wait2187;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2184\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 10;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0001" & \$v2184\&X"000000000";
                    state_var2250 <= pause_setI2185;
                  end if;
                when pause_setII2196 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2193\ := \$arr1646_ptr_take\;
                  if \$v2193\(0) = '1' then
                    state_var2250 <= q_wait2192;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2189\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 9;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0110" & \$v2189\&X"000000000";
                    state_var2250 <= pause_setI2190;
                  end if;
                when pause_setII2202 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2198\ := \$arr1646_ptr_take\;
                  if \$v2198\(0) = '1' then
                    state_var2250 <= q_wait2197;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2194\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 8;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2194\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2195;
                  end if;
                when pause_setII2207 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2204\ := \$arr1646_ptr_take\;
                  if \$v2204\(0) = '1' then
                    state_var2250 <= q_wait2203;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2199\ := eclat_unit;
                    \$v2200\ := "0010" & \$v2199\&"000"& X"000000000000000";
                    \$arr1646_ptr_write\ <= 7;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2200\;
                    state_var2250 <= pause_setI2201;
                  end if;
                when pause_setII2212 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2209\ := \$arr1646_ptr_take\;
                  if \$v2209\(0) = '1' then
                    state_var2250 <= q_wait2208;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2205\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 6;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2205\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2206;
                  end if;
                when pause_setII2219 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2214\ := \$arr1646_ptr_take\;
                  if \$v2214\(0) = '1' then
                    state_var2250 <= q_wait2213;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2210\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 5;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2210\&X"000000000";
                    state_var2250 <= pause_setI2211;
                  end if;
                when pause_setII2224 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2221\ := \$arr1646_ptr_take\;
                  if \$v2221\(0) = '1' then
                    state_var2250 <= q_wait2220;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2215\ := eclat_unit;
                    \$v2216\ := "0000" & \$v2215\;
                    \$v2217\ := "0011" & \$v2216\&"000"& X"00000000000000";
                    \$arr1646_ptr_write\ <= 4;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2217\;
                    state_var2250 <= pause_setI2218;
                  end if;
                when pause_setII2229 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2226\ := \$arr1646_ptr_take\;
                  if \$v2226\(0) = '1' then
                    state_var2250 <= q_wait2225;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2222\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 3;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2222\&X"000000000";
                    state_var2250 <= pause_setI2223;
                  end if;
                when pause_setII2234 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2231\ := \$arr1646_ptr_take\;
                  if \$v2231\(0) = '1' then
                    state_var2250 <= q_wait2230;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2227\ := "00000000000000000000000000000001";
                    \$arr1646_ptr_write\ <= 2;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2227\&X"000000000";
                    state_var2250 <= pause_setI2228;
                  end if;
                when pause_setII2239 =>
                  \$arr1646_ptr_take\(0) := '0';
                  \$v2236\ := \$arr1646_ptr_take\;
                  if \$v2236\(0) = '1' then
                    state_var2250 <= q_wait2235;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2232\ := "00000000000000000000000000001001";
                    \$arr1646_ptr_write\ <= 1;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1010" & \$v2232\&X"000000000";
                    state_var2250 <= pause_setI2233;
                  end if;
                when q_wait2116 =>
                  \$v2117\ := \$arr1643_ptr_take\;
                  if \$v2117\(0) = '1' then
                    state_var2250 <= q_wait2116;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr_write\ <= to_integer(unsigned(\$400_copy_args_to_heap518_arg\(64 to 95)));
                    \$arr1643_write_request\ <= '1';
                    \$arr1643_write\ <= \$593\;
                    state_var2250 <= pause_setI2114;
                  end if;
                when q_wait2120 =>
                  \$v2121\ := \$arr1644_ptr_take\;
                  if \$v2121\(0) = '1' then
                    state_var2250 <= q_wait2120;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$400_copy_args_to_heap518_arg\(32 to 63) & \$400_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var2250 <= pause_getI2118;
                  end if;
                when q_wait2130 =>
                  \$v2131\ := \$arr1644_ptr_take\;
                  if \$v2131\(0) = '1' then
                    state_var2250 <= q_wait2130;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$402_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$402_div543_arg\(0 to 31))));
                    state_var2250 <= pause_getI2128;
                  end if;
                when q_wait2138 =>
                  \$v2139\ := \$arr1644_ptr_take\;
                  if \$v2139\(0) = '1' then
                    state_var2250 <= q_wait2138;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$403_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$403_mul544_arg\(0 to 31))));
                    state_var2250 <= pause_getI2136;
                  end if;
                when q_wait2146 =>
                  \$v2147\ := \$arr1644_ptr_take\;
                  if \$v2147\(0) = '1' then
                    state_var2250 <= q_wait2146;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$404_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$404_sub545_arg\(0 to 31))));
                    state_var2250 <= pause_getI2144;
                  end if;
                when q_wait2154 =>
                  \$v2155\ := \$arr1644_ptr_take\;
                  if \$v2155\(0) = '1' then
                    state_var2250 <= q_wait2154;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$405_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$405_add546_arg\(0 to 31))));
                    state_var2250 <= pause_getI2152;
                  end if;
                when q_wait2160 =>
                  \$v2161\ := \$arr1646_ptr_take\;
                  if \$v2161\(0) = '1' then
                    state_var2250 <= q_wait2160;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2157\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 15;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0111" & \$v2157\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2158;
                  end if;
                when q_wait2165 =>
                  \$v2166\ := \$arr1646_ptr_take\;
                  if \$v2166\(0) = '1' then
                    state_var2250 <= q_wait2165;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2162\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 14;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2162\&X"000000000";
                    state_var2250 <= pause_setI2163;
                  end if;
                when q_wait2170 =>
                  \$v2171\ := \$arr1646_ptr_take\;
                  if \$v2171\(0) = '1' then
                    state_var2250 <= q_wait2170;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2167\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 13;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0010" & \$v2167\&X"000000000";
                    state_var2250 <= pause_setI2168;
                  end if;
                when q_wait2176 =>
                  \$v2177\ := \$arr1646_ptr_take\;
                  if \$v2177\(0) = '1' then
                    state_var2250 <= q_wait2176;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2172\ := "00000000000000000000000000000001";
                    \$v2173\ := "0001" & \$v2172\&X"00000000";
                    \$arr1646_ptr_write\ <= 12;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2173\;
                    state_var2250 <= pause_setI2174;
                  end if;
                when q_wait2182 =>
                  \$v2183\ := \$arr1646_ptr_take\;
                  if \$v2183\(0) = '1' then
                    state_var2250 <= q_wait2182;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2178\ := "00000000000000000000000000000010";
                    \$v2179\ := "0001" & \$v2178\&X"00000000";
                    \$arr1646_ptr_write\ <= 11;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2179\;
                    state_var2250 <= pause_setI2180;
                  end if;
                when q_wait2187 =>
                  \$v2188\ := \$arr1646_ptr_take\;
                  if \$v2188\(0) = '1' then
                    state_var2250 <= q_wait2187;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2184\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 10;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0001" & \$v2184\&X"000000000";
                    state_var2250 <= pause_setI2185;
                  end if;
                when q_wait2192 =>
                  \$v2193\ := \$arr1646_ptr_take\;
                  if \$v2193\(0) = '1' then
                    state_var2250 <= q_wait2192;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2189\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 9;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0110" & \$v2189\&X"000000000";
                    state_var2250 <= pause_setI2190;
                  end if;
                when q_wait2197 =>
                  \$v2198\ := \$arr1646_ptr_take\;
                  if \$v2198\(0) = '1' then
                    state_var2250 <= q_wait2197;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2194\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 8;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2194\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2195;
                  end if;
                when q_wait2203 =>
                  \$v2204\ := \$arr1646_ptr_take\;
                  if \$v2204\(0) = '1' then
                    state_var2250 <= q_wait2203;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2199\ := eclat_unit;
                    \$v2200\ := "0010" & \$v2199\&"000"& X"000000000000000";
                    \$arr1646_ptr_write\ <= 7;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2200\;
                    state_var2250 <= pause_setI2201;
                  end if;
                when q_wait2208 =>
                  \$v2209\ := \$arr1646_ptr_take\;
                  if \$v2209\(0) = '1' then
                    state_var2250 <= q_wait2208;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2205\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 6;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1001" & \$v2205\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2206;
                  end if;
                when q_wait2213 =>
                  \$v2214\ := \$arr1646_ptr_take\;
                  if \$v2214\(0) = '1' then
                    state_var2250 <= q_wait2213;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2210\ := "00000000000000000000000000000010";
                    \$arr1646_ptr_write\ <= 5;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1000" & \$v2210\&X"000000000";
                    state_var2250 <= pause_setI2211;
                  end if;
                when q_wait2220 =>
                  \$v2221\ := \$arr1646_ptr_take\;
                  if \$v2221\(0) = '1' then
                    state_var2250 <= q_wait2220;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2215\ := eclat_unit;
                    \$v2216\ := "0000" & \$v2215\;
                    \$v2217\ := "0011" & \$v2216\&"000"& X"00000000000000";
                    \$arr1646_ptr_write\ <= 4;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0101" & \$v2217\;
                    state_var2250 <= pause_setI2218;
                  end if;
                when q_wait2225 =>
                  \$v2226\ := \$arr1646_ptr_take\;
                  if \$v2226\(0) = '1' then
                    state_var2250 <= q_wait2225;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2222\ := "00000000000000000000000000000000";
                    \$arr1646_ptr_write\ <= 3;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2222\&X"000000000";
                    state_var2250 <= pause_setI2223;
                  end if;
                when q_wait2230 =>
                  \$v2231\ := \$arr1646_ptr_take\;
                  if \$v2231\(0) = '1' then
                    state_var2250 <= q_wait2230;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2227\ := "00000000000000000000000000000001";
                    \$arr1646_ptr_write\ <= 2;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0100" & \$v2227\&X"000000000";
                    state_var2250 <= pause_setI2228;
                  end if;
                when q_wait2235 =>
                  \$v2236\ := \$arr1646_ptr_take\;
                  if \$v2236\(0) = '1' then
                    state_var2250 <= q_wait2235;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2232\ := "00000000000000000000000000001001";
                    \$arr1646_ptr_write\ <= 1;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "1010" & \$v2232\&X"000000000";
                    state_var2250 <= pause_setI2233;
                  end if;
                when q_wait2240 =>
                  \$v2241\ := \$arr1646_ptr_take\;
                  if \$v2241\(0) = '1' then
                    state_var2250 <= q_wait2240;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2237\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 0;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0000" & \$v2237\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2238;
                  end if;
                when compute2113 =>
                  rdy2112 := eclat_false;
                  \$v2241\ := \$arr1646_ptr_take\;
                  if \$v2241\(0) = '1' then
                    state_var2250 <= q_wait2240;
                  else
                    \$arr1646_ptr_take\(0) := '1';
                    \$v2237\ := eclat_unit;
                    \$arr1646_ptr_write\ <= 0;
                    \$arr1646_write_request\ <= '1';
                    \$arr1646_write\ <= "0000" & \$v2237\&"000"& X"0000000000000000";
                    state_var2250 <= pause_setI2238;
                  end if;
                end case;
                \$v2243\ := eclat_not(rdy2112);
                if \$v2243\(0) = '1' then
                  result2111 := eclat_unit;
                end if;
                \$397\ := result2111 & rdy2112;
                result2108 := ""&\$397\(1);
                rdy2109 := eclat_true;
                state_var2249 <= compute2110;
              end if;
            end case;
            \$v2246\ := eclat_not(rdy2109);
            if \$v2246\(0) = '1' then
              result2108 := eclat_false;
            end if;
            \$395\ := result2108;
            \$134_is_loaded\ := result2108;
            case state_var2248 is
            when compute2105 =>
              rdy2104 := eclat_false;
              result2103 := eclat_if(\$134_is_loaded\ & eclat_add(\$393\ & "00000000000000000000000000000001") & \$393\);
              rdy2104 := eclat_true;
              state_var2248 <= compute2105;
            end case;
            \$v2107\ := eclat_not(rdy2104);
            if \$v2107\(0) = '1' then
              result2103 := "00000000000000000000000000000000";
            end if;
            \$393\ := result2103;
            \$135_cy\ := result2103;
            case state_var2247 is
            when \$117_forever5471614\ =>
              state_var2247 <= \$117_forever5471614\;
            when \$117_forever5471621\ =>
              state_var2247 <= \$117_forever5471614\;
            when \$117_forever5471622\ =>
              state_var2247 <= \$117_forever5471614\;
            when \$117_forever5471623\ =>
              state_var2247 <= \$117_forever5471614\;
            when \$117_forever5471624\ =>
              state_var2247 <= \$117_forever5471614\;
            when \$120_forever5481613\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481625\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481626\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481627\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481628\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481629\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481630\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481631\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481632\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481633\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481634\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$120_forever5481635\ =>
              state_var2247 <= \$120_forever5481613\;
            when \$143_copy_args_to_heap518\ =>
              \$v1706\ := eclat_eq(\$143_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1706\(0) = '1' then
                \$143_copy_args_to_heap518_result\ := \$143_copy_args_to_heap518_arg\(32 to 63);
                \$v1751\ := \$arr1647_ptr_take\;
                if \$v1751\(0) = '1' then
                  state_var2247 <= q_wait1750;
                else
                  \$arr1647_ptr_take\(0) := '1';
                  \$arr1647_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(96 to 127)));
                  \$arr1647_write_request\ <= '1';
                  \$arr1647_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127);
                  state_var2247 <= pause_setI1748;
                end if;
              else
                \$v1705\ := \$arr1644_ptr_take\;
                if \$v1705\(0) = '1' then
                  state_var2247 <= q_wait1704;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$143_copy_args_to_heap518_arg\(32 to 63) & \$143_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1702;
                end if;
              end if;
            when \$144_pow542\ =>
              \$v1707\ := eclat_eq(\$144_pow542_arg\(32 to 63) & "00000000000000000000000000000000");
              if \$v1707\(0) = '1' then
                \$144_pow542_result\ := \$144_pow542_arg\(64 to 95);
                resultat := \$144_pow542_result\;
                \$v1847\ := \$arr1644_ptr_take\;
                if \$v1847\(0) = '1' then
                  state_var2247 <= q_wait1846;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1844;
                end if;
              else
                \$144_pow542_arg\ := \$144_pow542_arg\(0 to 31) & eclat_sub(\$144_pow542_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$144_pow542_arg\(64 to 95) & \$144_pow542_arg\(0 to 31));
                state_var2247 <= \$144_pow542\;
              end if;
            when \$145_div543\ =>
              \$v1716\ := eclat_eq(\$145_div543_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1716\(0) = '1' then
                \$145_div543_result\ := \$145_div543_arg\(32 to 63);
                resultat := \$145_div543_result\;
                \$v1866\ := \$arr1644_ptr_take\;
                if \$v1866\(0) = '1' then
                  state_var2247 <= q_wait1865;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1863;
                end if;
              else
                \$v1715\ := \$arr1644_ptr_take\;
                if \$v1715\(0) = '1' then
                  state_var2247 <= q_wait1714;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$145_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$145_div543_arg\(0 to 31))));
                  state_var2247 <= pause_getI1712;
                end if;
              end if;
            when \$146_mul544\ =>
              \$v1724\ := eclat_eq(\$146_mul544_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1724\(0) = '1' then
                \$146_mul544_result\ := \$146_mul544_arg\(32 to 63);
                resultat := \$146_mul544_result\;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1911\ := \$arr1644_ptr_take\;
                if \$v1911\(0) = '1' then
                  state_var2247 <= q_wait1910;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1908;
                end if;
              else
                \$v1723\ := \$arr1644_ptr_take\;
                if \$v1723\(0) = '1' then
                  state_var2247 <= q_wait1722;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_mul544_arg\(0 to 31))));
                  state_var2247 <= pause_getI1720;
                end if;
              end if;
            when \$147_sub545\ =>
              \$v1732\ := eclat_eq(\$147_sub545_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1732\(0) = '1' then
                \$147_sub545_result\ := \$147_sub545_arg\(32 to 63);
                resultat := \$147_sub545_result\;
                \$v1916\ := \$arr1644_ptr_take\;
                if \$v1916\(0) = '1' then
                  state_var2247 <= q_wait1915;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1912\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & \$v1912\&X"00000000";
                  state_var2247 <= pause_setI1913;
                end if;
              else
                \$v1731\ := \$arr1644_ptr_take\;
                if \$v1731\(0) = '1' then
                  state_var2247 <= q_wait1730;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_sub545_arg\(0 to 31))));
                  state_var2247 <= pause_getI1728;
                end if;
              end if;
            when \$148_add546\ =>
              \$v1740\ := eclat_eq(\$148_add546_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1740\(0) = '1' then
                \$148_add546_result\ := \$148_add546_arg\(32 to 63);
                resultat := \$148_add546_result\;
                \$v1961\ := \$arr1644_ptr_take\;
                if \$v1961\(0) = '1' then
                  state_var2247 <= q_wait1960;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1958;
                end if;
              else
                \$v1739\ := \$arr1644_ptr_take\;
                if \$v1739\(0) = '1' then
                  state_var2247 <= q_wait1738;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_add546_arg\(0 to 31))));
                  state_var2247 <= pause_getI1736;
                end if;
              end if;
            when \$149_vm_run_code521\ =>
              \$v2099\ := ""&\$149_vm_run_code521_arg\(294);
              if \$v2099\(0) = '1' then
                eclat_print_string(of_string("[sp:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(0 to 31));
                
                eclat_print_string(of_string("|env:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(32 to 63));
                
                eclat_print_string(of_string("|pc:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(64 to 95));
                
                eclat_print_string(of_string("|fp:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(96 to 127));
                
                eclat_print_string(of_string("]"));
                
                eclat_print_string(of_string("|gp:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(128 to 159));
                
                eclat_print_string(of_string("|hp:"));
                
                eclat_print_int(\$149_vm_run_code521_arg\(128 to 159));
                
                eclat_print_newline(eclat_unit);
                
                \$v2098\ := \$arr1646_ptr_take\;
                if \$v2098\(0) = '1' then
                  state_var2247 <= q_wait2097;
                else
                  \$arr1646_ptr_take\(0) := '1';
                  \$arr1646_ptr\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(64 to 95)));
                  state_var2247 <= pause_getI2095;
                end if;
              else
                \$v2098\ := \$arr1646_ptr_take\;
                if \$v2098\(0) = '1' then
                  state_var2247 <= q_wait2097;
                else
                  \$arr1646_ptr_take\(0) := '1';
                  \$arr1646_ptr\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(64 to 95)));
                  state_var2247 <= pause_getI2095;
                end if;
              end if;
            when \$208_forever5471620\ =>
              state_var2247 <= \$212_forever5471614\;
            when \$212_forever5471614\ =>
              state_var2247 <= \$212_forever5471614\;
            when \$258_forever5481619\ =>
              state_var2247 <= \$262_forever5481613\;
            when \$262_forever5481613\ =>
              state_var2247 <= \$262_forever5481613\;
            when \$287_forever5481618\ =>
              state_var2247 <= \$291_forever5481613\;
            when \$291_forever5481613\ =>
              state_var2247 <= \$291_forever5481613\;
            when \$316_forever5481617\ =>
              state_var2247 <= \$320_forever5481613\;
            when \$320_forever5481613\ =>
              state_var2247 <= \$320_forever5481613\;
            when \$344_forever5481615\ =>
              state_var2247 <= \$348_forever5481613\;
            when \$348_forever5481613\ =>
              state_var2247 <= \$348_forever5481613\;
            when \$357_forever5481616\ =>
              state_var2247 <= \$361_forever5481613\;
            when \$361_forever5481613\ =>
              state_var2247 <= \$361_forever5481613\;
            when pause_getI1702 =>
              state_var2247 <= pause_getII1703;
            when pause_getI1712 =>
              state_var2247 <= pause_getII1713;
            when pause_getI1720 =>
              state_var2247 <= pause_getII1721;
            when pause_getI1728 =>
              state_var2247 <= pause_getII1729;
            when pause_getI1736 =>
              state_var2247 <= pause_getII1737;
            when pause_getI1774 =>
              state_var2247 <= pause_getII1775;
            when pause_getI1778 =>
              state_var2247 <= pause_getII1779;
            when pause_getI1803 =>
              state_var2247 <= pause_getII1804;
            when pause_getI1814 =>
              state_var2247 <= pause_getII1815;
            when pause_getI1825 =>
              state_var2247 <= pause_getII1826;
            when pause_getI1832 =>
              state_var2247 <= pause_getII1833;
            when pause_getI1839 =>
              state_var2247 <= pause_getII1840;
            when pause_getI1851 =>
              state_var2247 <= pause_getII1852;
            when pause_getI1858 =>
              state_var2247 <= pause_getII1859;
            when pause_getI1870 =>
              state_var2247 <= pause_getII1871;
            when pause_getI1886 =>
              state_var2247 <= pause_getII1887;
            when pause_getI1897 =>
              state_var2247 <= pause_getII1898;
            when pause_getI1908 =>
              state_var2247 <= pause_getII1909;
            when pause_getI1924 =>
              state_var2247 <= pause_getII1925;
            when pause_getI1935 =>
              state_var2247 <= pause_getII1936;
            when pause_getI1946 =>
              state_var2247 <= pause_getII1947;
            when pause_getI1953 =>
              state_var2247 <= pause_getII1954;
            when pause_getI1969 =>
              state_var2247 <= pause_getII1970;
            when pause_getI1980 =>
              state_var2247 <= pause_getII1981;
            when pause_getI1991 =>
              state_var2247 <= pause_getII1992;
            when pause_getI1999 =>
              state_var2247 <= pause_getII2000;
            when pause_getI2012 =>
              state_var2247 <= pause_getII2013;
            when pause_getI2016 =>
              state_var2247 <= pause_getII2017;
            when pause_getI2023 =>
              state_var2247 <= pause_getII2024;
            when pause_getI2030 =>
              state_var2247 <= pause_getII2031;
            when pause_getI2038 =>
              state_var2247 <= pause_getII2039;
            when pause_getI2046 =>
              state_var2247 <= pause_getII2047;
            when pause_getI2057 =>
              state_var2247 <= pause_getII2058;
            when pause_getI2065 =>
              state_var2247 <= pause_getII2066;
            when pause_getI2073 =>
              state_var2247 <= pause_getII2074;
            when pause_getI2084 =>
              state_var2247 <= pause_getII2085;
            when pause_getI2095 =>
              state_var2247 <= pause_getII2096;
            when pause_getII1703 =>
              \$arr1644_ptr_take\(0) := '0';
              \$389\ := \$arr1644_value\;
              \$v1701\ := \$arr1643_ptr_take\;
              if \$v1701\(0) = '1' then
                state_var2247 <= q_wait1700;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(\$143_copy_args_to_heap518_arg\(64 to 95)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= \$389\;
                state_var2247 <= pause_setI1698;
              end if;
            when pause_getII1713 =>
              \$arr1644_ptr_take\(0) := '0';
              \$352\ := \$arr1644_value\;
              \$v1710\ := \$352\;
              \$v1711\ := \$v1710\(0 to 3);
              \$v1709\ := \$v1710\(4 to 67);
              case \$v1711\ is
              when "0001" =>
                \$353_a\ := \$v1709\(0 to 31);
                \$335_divisor\ := \$353_a\;
                \$v1708\ := eclat_eq(\$335_divisor\ & "00000000000000000000000000000000");
                if \$v1708\(0) = '1' then
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("Division par zero"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2247 <= \$344_forever5481615\;
                else
                  \$145_div543_arg\ := eclat_sub(\$145_div543_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$145_div543_arg\(32 to 63) & \$335_divisor\) & \$145_div543_arg\(64 to 95);
                  state_var2247 <= \$145_div543\;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$357_forever5481616\;
              end case;
            when pause_getII1721 =>
              \$arr1644_ptr_take\(0) := '0';
              \$306_v\ := \$arr1644_value\;
              \$v1718\ := \$306_v\;
              \$v1719\ := \$v1718\(0 to 3);
              \$v1717\ := \$v1718\(4 to 67);
              case \$v1719\ is
              when "0001" =>
                \$312_a\ := \$v1717\(0 to 31);
                \$307_int_value\ := \$312_a\;
                \$146_mul544_arg\ := eclat_sub(\$146_mul544_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$146_mul544_arg\(32 to 63) & \$307_int_value\) & \$146_mul544_arg\(64 to 95);
                state_var2247 <= \$146_mul544\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$316_forever5481617\;
              end case;
            when pause_getII1729 =>
              \$arr1644_ptr_take\(0) := '0';
              \$277_v\ := \$arr1644_value\;
              \$v1726\ := \$277_v\;
              \$v1727\ := \$v1726\(0 to 3);
              \$v1725\ := \$v1726\(4 to 67);
              case \$v1727\ is
              when "0001" =>
                \$283_a\ := \$v1725\(0 to 31);
                \$278_int_value\ := \$283_a\;
                \$147_sub545_arg\ := eclat_sub(\$147_sub545_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$147_sub545_arg\(32 to 63) & \$278_int_value\) & \$147_sub545_arg\(64 to 95);
                state_var2247 <= \$147_sub545\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$287_forever5481618\;
              end case;
            when pause_getII1737 =>
              \$arr1644_ptr_take\(0) := '0';
              \$248_v\ := \$arr1644_value\;
              \$v1734\ := \$248_v\;
              \$v1735\ := \$v1734\(0 to 3);
              \$v1733\ := \$v1734\(4 to 67);
              case \$v1735\ is
              when "0001" =>
                \$254_a\ := \$v1733\(0 to 31);
                \$249_int_value\ := \$254_a\;
                \$148_add546_arg\ := eclat_sub(\$148_add546_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$148_add546_arg\(32 to 63) & \$249_int_value\) & \$148_add546_arg\(64 to 95);
                state_var2247 <= \$148_add546\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur dans ADD, c'est pas un entier "));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$258_forever5481619\;
              end case;
            when pause_getII1775 =>
              \$arr1644_ptr_take\(0) := '0';
              second_value := \$arr1644_value\;
              \$v1772\ := first_value;
              \$v1773\ := \$v1772\(0 to 3);
              \$v1762\ := \$v1772\(4 to 67);
              case \$v1773\ is
              when "0010" =>
                \$v1764\ := second_value;
                \$v1765\ := \$v1764\(0 to 3);
                \$v1763\ := \$v1764\(4 to 67);
                case \$v1765\ is
                when "0010" =>
                  res := eclat_true;
                  \$v1761\ := \$arr1644_ptr_take\;
                  if \$v1761\(0) = '1' then
                    state_var2247 <= q_wait1760;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1758;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2247 <= \$117_forever5471622\;
                end case;
              when "0000" =>
                \$98_a1\ := \$v1762\(0 to 0);
                \$v1767\ := second_value;
                \$v1768\ := \$v1767\(0 to 3);
                \$v1766\ := \$v1767\(4 to 67);
                case \$v1768\ is
                when "0000" =>
                  b2 := \$v1766\(0 to 0);
                  res := eclat_if(\$98_a1\ & eclat_if(b2 & eclat_true & eclat_false) & 
                         eclat_if(b2 & eclat_false & eclat_true));
                  \$v1761\ := \$arr1644_ptr_take\;
                  if \$v1761\(0) = '1' then
                    state_var2247 <= q_wait1760;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1758;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2247 <= \$117_forever5471623\;
                end case;
              when "0001" =>
                \$99_a\ := \$v1762\(0 to 31);
                \$v1770\ := second_value;
                \$v1771\ := \$v1770\(0 to 3);
                \$v1769\ := \$v1770\(4 to 67);
                case \$v1771\ is
                when "0001" =>
                  b := \$v1769\(0 to 31);
                  res := eclat_eq(\$99_a\ & b);
                  \$v1761\ := \$arr1644_ptr_take\;
                  if \$v1761\(0) = '1' then
                    state_var2247 <= q_wait1760;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1758;
                  end if;
                when others =>
                  eclat_print_string(of_string("types incompatibles\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var2247 <= \$117_forever5471624\;
                end case;
              when others =>
                eclat_print_string(of_string("il n'y a pas d'égalité possible \n"));
                
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$117_forever5471621\;
              end case;
            when pause_getII1779 =>
              \$arr1644_ptr_take\(0) := '0';
              first_value := \$arr1644_value\;
              \$v1777\ := \$arr1644_ptr_take\;
              if \$v1777\(0) = '1' then
                state_var2247 <= q_wait1776;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2247 <= pause_getI1774;
              end if;
            when pause_getII1804 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v56\ := \$arr1644_value\;
              \$v1801\ := \$v56\;
              \$v1802\ := \$v1801\(0 to 3);
              \$v1796\ := \$v1801\(4 to 67);
              case \$v1802\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1795\ := \$arr1644_ptr_take\;
                if \$v1795\(0) = '1' then
                  state_var2247 <= q_wait1794;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1791\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                  state_var2247 <= pause_setI1792;
                end if;
              when "0011" =>
                \$113_p\ := \$v1796\(0 to 4);
                \$v1798\ := \$113_p\;
                \$v1799\ := \$v1798\(0 to 3);
                \$v1797\ := ""&\$v1798\(4);
                case \$v1799\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1795\ := \$arr1644_ptr_take\;
                if \$v1795\(0) = '1' then
                  state_var2247 <= q_wait1794;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1791\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                  state_var2247 <= pause_setI1792;
                end if;
              when "0001" =>
                \$114_n\ := \$v1796\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v1795\ := \$arr1644_ptr_take\;
                if \$v1795\(0) = '1' then
                  state_var2247 <= q_wait1794;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v1791\ := eclat_gt(fst_operand & scd_operand);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                  state_var2247 <= pause_setI1792;
                end if;
              when "0000" =>
                \$115_b\ := \$v1796\(0 to 0);
                \$v1800\ := \$115_b\;
                if \$v1800\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1795\ := \$arr1644_ptr_take\;
                  if \$v1795\(0) = '1' then
                    state_var2247 <= q_wait1794;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$v1791\ := eclat_gt(fst_operand & scd_operand);
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                    state_var2247 <= pause_setI1792;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1815 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v53\ := \$arr1644_value\;
              \$v1812\ := \$v53\;
              \$v1813\ := \$v1812\(0 to 3);
              \$v1807\ := \$v1812\(4 to 67);
              case \$v1813\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1806\ := \$arr1644_ptr_take\;
                if \$v1806\(0) = '1' then
                  state_var2247 <= q_wait1805;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1803;
                end if;
              when "0011" =>
                \$113_p\ := \$v1807\(0 to 4);
                \$v1809\ := \$113_p\;
                \$v1810\ := \$v1809\(0 to 3);
                \$v1808\ := ""&\$v1809\(4);
                case \$v1810\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1806\ := \$arr1644_ptr_take\;
                if \$v1806\(0) = '1' then
                  state_var2247 <= q_wait1805;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1803;
                end if;
              when "0001" =>
                \$114_n\ := \$v1807\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1806\ := \$arr1644_ptr_take\;
                if \$v1806\(0) = '1' then
                  state_var2247 <= q_wait1805;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1803;
                end if;
              when "0000" =>
                \$115_b\ := \$v1807\(0 to 0);
                \$v1811\ := \$115_b\;
                if \$v1811\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1806\ := \$arr1644_ptr_take\;
                  if \$v1806\(0) = '1' then
                    state_var2247 <= q_wait1805;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1803;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1826 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v50\ := \$arr1644_value\;
              \$v1823\ := \$v50\;
              \$v1824\ := \$v1823\(0 to 3);
              \$v1818\ := \$v1823\(4 to 67);
              case \$v1824\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2247 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2247 <= pause_getI1814;
                end if;
              when "0011" =>
                \$113_p\ := \$v1818\(0 to 4);
                \$v1820\ := \$113_p\;
                \$v1821\ := \$v1820\(0 to 3);
                \$v1819\ := ""&\$v1820\(4);
                case \$v1821\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2247 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2247 <= pause_getI1814;
                end if;
              when "0001" =>
                \$114_n\ := \$v1818\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1817\ := \$arr1644_ptr_take\;
                if \$v1817\(0) = '1' then
                  state_var2247 <= q_wait1816;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2247 <= pause_getI1814;
                end if;
              when "0000" =>
                \$115_b\ := \$v1818\(0 to 0);
                \$v1822\ := \$115_b\;
                if \$v1822\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1817\ := \$arr1644_ptr_take\;
                  if \$v1817\(0) = '1' then
                    state_var2247 <= q_wait1816;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                    state_var2247 <= pause_getI1814;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1833 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v47\ := \$arr1644_value\;
              \$v1830\ := \$v47\;
              \$v1831\ := \$v1830\(0 to 3);
              \$v1829\ := \$v1830\(4 to 67);
              case \$v1831\ is
              when "0001" =>
                a := \$v1829\(0 to 31);
                scd_operand := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1828\ := \$arr1644_ptr_take\;
                if \$v1828\(0) = '1' then
                  state_var2247 <= q_wait1827;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                  state_var2247 <= pause_getI1825;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481626\;
              end case;
            when pause_getII1840 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v45\ := \$arr1644_value\;
              \$v1837\ := \$v45\;
              \$v1838\ := \$v1837\(0 to 3);
              \$v1836\ := \$v1837\(4 to 67);
              case \$v1838\ is
              when "0001" =>
                a := \$v1836\(0 to 31);
                fst_operand := a;
                \$v1835\ := \$arr1644_ptr_take\;
                if \$v1835\(0) = '1' then
                  state_var2247 <= q_wait1834;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2247 <= pause_getI1832;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481627\;
              end case;
            when pause_getII1852 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v68\ := \$arr1644_value\;
              \$v1849\ := \$v68\;
              \$v1850\ := \$v1849\(0 to 3);
              \$v1848\ := \$v1849\(4 to 67);
              case \$v1850\ is
              when "0001" =>
                a := \$v1848\(0 to 31);
                exponent := a;
                \$144_pow542_arg\ := base & exponent & "00000000000000000000000000000001";
                state_var2247 <= \$144_pow542\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481629\;
              end case;
            when pause_getII1859 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v66\ := \$arr1644_value\;
              \$v1856\ := \$v66\;
              \$v1857\ := \$v1856\(0 to 3);
              \$v1855\ := \$v1856\(4 to 67);
              case \$v1857\ is
              when "0001" =>
                a := \$v1855\(0 to 31);
                base := a;
                \$v1854\ := \$arr1644_ptr_take\;
                if \$v1854\(0) = '1' then
                  state_var2247 <= q_wait1853;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                  state_var2247 <= pause_getI1851;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481630\;
              end case;
            when pause_getII1871 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v92\ := \$arr1644_value\;
              \$v1868\ := \$v92\;
              \$v1869\ := \$v1868\(0 to 3);
              \$v1867\ := \$v1868\(4 to 67);
              case \$v1869\ is
              when "0001" =>
                a := \$v1867\(0 to 31);
                debut := a;
                \$145_div543_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$145_div543\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481632\;
              end case;
            when pause_getII1887 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v124\ := \$arr1644_value\;
              \$v1884\ := \$v124\;
              \$v1885\ := \$v1884\(0 to 3);
              \$v1879\ := \$v1884\(4 to 67);
              case \$v1885\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1878\ := \$arr1644_ptr_take\;
                if \$v1878\(0) = '1' then
                  state_var2247 <= q_wait1877;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1875;
                end if;
              when "0011" =>
                \$113_p\ := \$v1879\(0 to 4);
                \$v1881\ := \$113_p\;
                \$v1882\ := \$v1881\(0 to 3);
                \$v1880\ := ""&\$v1881\(4);
                case \$v1882\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v1878\ := \$arr1644_ptr_take\;
                if \$v1878\(0) = '1' then
                  state_var2247 <= q_wait1877;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1875;
                end if;
              when "0001" =>
                \$114_n\ := \$v1879\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v1878\ := \$arr1644_ptr_take\;
                if \$v1878\(0) = '1' then
                  state_var2247 <= q_wait1877;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0001" & resultat&X"00000000";
                  state_var2247 <= pause_setI1875;
                end if;
              when "0000" =>
                \$115_b\ := \$v1879\(0 to 0);
                \$v1883\ := \$115_b\;
                if \$v1883\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v1878\ := \$arr1644_ptr_take\;
                  if \$v1878\(0) = '1' then
                    state_var2247 <= q_wait1877;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    \$arr1644_write_request\ <= '1';
                    \$arr1644_write\ <= "0001" & resultat&X"00000000";
                    state_var2247 <= pause_setI1875;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1898 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v117\ := \$arr1644_value\;
              \$v1895\ := \$v117\;
              \$v1896\ := \$v1895\(0 to 3);
              \$v1890\ := \$v1895\(4 to 67);
              case \$v1896\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1889\ := \$arr1644_ptr_take\;
                if \$v1889\(0) = '1' then
                  state_var2247 <= q_wait1888;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1886;
                end if;
              when "0011" =>
                \$113_p\ := \$v1890\(0 to 4);
                \$v1892\ := \$113_p\;
                \$v1893\ := \$v1892\(0 to 3);
                \$v1891\ := ""&\$v1892\(4);
                case \$v1893\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1889\ := \$arr1644_ptr_take\;
                if \$v1889\(0) = '1' then
                  state_var2247 <= q_wait1888;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1886;
                end if;
              when "0001" =>
                \$114_n\ := \$v1890\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1889\ := \$arr1644_ptr_take\;
                if \$v1889\(0) = '1' then
                  state_var2247 <= q_wait1888;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1886;
                end if;
              when "0000" =>
                \$115_b\ := \$v1890\(0 to 0);
                \$v1894\ := \$115_b\;
                if \$v1894\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1889\ := \$arr1644_ptr_take\;
                  if \$v1889\(0) = '1' then
                    state_var2247 <= q_wait1888;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1886;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1909 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v114\ := \$arr1644_value\;
              \$v1906\ := \$v114\;
              \$v1907\ := \$v1906\(0 to 3);
              \$v1901\ := \$v1906\(4 to 67);
              case \$v1907\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2247 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1897;
                end if;
              when "0011" =>
                \$113_p\ := \$v1901\(0 to 4);
                \$v1903\ := \$113_p\;
                \$v1904\ := \$v1903\(0 to 3);
                \$v1902\ := ""&\$v1903\(4);
                case \$v1904\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2247 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1897;
                end if;
              when "0001" =>
                \$114_n\ := \$v1901\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1900\ := \$arr1644_ptr_take\;
                if \$v1900\(0) = '1' then
                  state_var2247 <= q_wait1899;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1897;
                end if;
              when "0000" =>
                \$115_b\ := \$v1901\(0 to 0);
                \$v1905\ := \$115_b\;
                if \$v1905\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1900\ := \$arr1644_ptr_take\;
                  if \$v1900\(0) = '1' then
                    state_var2247 <= q_wait1899;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1897;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1925 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v159\ := \$arr1644_value\;
              \$v1922\ := \$v159\;
              \$v1923\ := \$v1922\(0 to 3);
              \$v1917\ := \$v1922\(4 to 67);
              case \$v1923\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$147_sub545\;
              when "0011" =>
                \$113_p\ := \$v1917\(0 to 4);
                \$v1919\ := \$113_p\;
                \$v1920\ := \$v1919\(0 to 3);
                \$v1918\ := ""&\$v1919\(4);
                case \$v1920\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$147_sub545\;
              when "0001" =>
                \$114_n\ := \$v1917\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$147_sub545\;
              when "0000" =>
                \$115_b\ := \$v1917\(0 to 0);
                \$v1921\ := \$115_b\;
                if \$v1921\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$147_sub545_arg\ := eclat_sub(\$192_n\ & "00000000000000000000000000000001") & debut & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$147_sub545\;
                end if;
              when others =>
                
              end case;
            when pause_getII1936 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v152\ := \$arr1644_value\;
              \$v1933\ := \$v152\;
              \$v1934\ := \$v1933\(0 to 3);
              \$v1928\ := \$v1933\(4 to 67);
              case \$v1934\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1927\ := \$arr1644_ptr_take\;
                if \$v1927\(0) = '1' then
                  state_var2247 <= q_wait1926;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1924;
                end if;
              when "0011" =>
                \$113_p\ := \$v1928\(0 to 4);
                \$v1930\ := \$113_p\;
                \$v1931\ := \$v1930\(0 to 3);
                \$v1929\ := ""&\$v1930\(4);
                case \$v1931\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1927\ := \$arr1644_ptr_take\;
                if \$v1927\(0) = '1' then
                  state_var2247 <= q_wait1926;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1924;
                end if;
              when "0001" =>
                \$114_n\ := \$v1928\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1927\ := \$arr1644_ptr_take\;
                if \$v1927\(0) = '1' then
                  state_var2247 <= q_wait1926;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1924;
                end if;
              when "0000" =>
                \$115_b\ := \$v1928\(0 to 0);
                \$v1932\ := \$115_b\;
                if \$v1932\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1927\ := \$arr1644_ptr_take\;
                  if \$v1927\(0) = '1' then
                    state_var2247 <= q_wait1926;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1924;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1947 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v149\ := \$arr1644_value\;
              \$v1944\ := \$v149\;
              \$v1945\ := \$v1944\(0 to 3);
              \$v1939\ := \$v1944\(4 to 67);
              case \$v1945\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1938\ := \$arr1644_ptr_take\;
                if \$v1938\(0) = '1' then
                  state_var2247 <= q_wait1937;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1935;
                end if;
              when "0011" =>
                \$113_p\ := \$v1939\(0 to 4);
                \$v1941\ := \$113_p\;
                \$v1942\ := \$v1941\(0 to 3);
                \$v1940\ := ""&\$v1941\(4);
                case \$v1942\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1938\ := \$arr1644_ptr_take\;
                if \$v1938\(0) = '1' then
                  state_var2247 <= q_wait1937;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1935;
                end if;
              when "0001" =>
                \$114_n\ := \$v1939\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1938\ := \$arr1644_ptr_take\;
                if \$v1938\(0) = '1' then
                  state_var2247 <= q_wait1937;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1935;
                end if;
              when "0000" =>
                \$115_b\ := \$v1939\(0 to 0);
                \$v1943\ := \$115_b\;
                if \$v1943\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1938\ := \$arr1644_ptr_take\;
                  if \$v1938\(0) = '1' then
                    state_var2247 <= q_wait1937;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1935;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1954 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v142\ := \$arr1644_value\;
              \$v1951\ := \$v142\;
              \$v1952\ := \$v1951\(0 to 3);
              \$v1950\ := \$v1951\(4 to 67);
              case \$v1952\ is
              when "0001" =>
                a := \$v1950\(0 to 31);
                debut := a;
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1949\ := \$arr1644_ptr_take\;
                if \$v1949\(0) = '1' then
                  state_var2247 <= q_wait1948;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1946;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("erreur"));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$120_forever5481634\;
              end case;
            when pause_getII1970 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v194\ := \$arr1644_value\;
              \$v1967\ := \$v194\;
              \$v1968\ := \$v1967\(0 to 3);
              \$v1962\ := \$v1967\(4 to 67);
              case \$v1968\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$148_add546\;
              when "0011" =>
                \$113_p\ := \$v1962\(0 to 4);
                \$v1964\ := \$113_p\;
                \$v1965\ := \$v1964\(0 to 3);
                \$v1963\ := ""&\$v1964\(4);
                case \$v1965\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$148_add546\;
              when "0001" =>
                \$114_n\ := \$v1962\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                state_var2247 <= \$148_add546\;
              when "0000" =>
                \$115_b\ := \$v1962\(0 to 0);
                \$v1966\ := \$115_b\;
                if \$v1966\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$148_add546_arg\ := \$192_n\ & "00000000000000000000000000000000" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$148_add546\;
                end if;
              when others =>
                
              end case;
            when pause_getII1981 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v187\ := \$arr1644_value\;
              \$v1978\ := \$v187\;
              \$v1979\ := \$v1978\(0 to 3);
              \$v1973\ := \$v1978\(4 to 67);
              case \$v1979\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1972\ := \$arr1644_ptr_take\;
                if \$v1972\(0) = '1' then
                  state_var2247 <= q_wait1971;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1969;
                end if;
              when "0011" =>
                \$113_p\ := \$v1973\(0 to 4);
                \$v1975\ := \$113_p\;
                \$v1976\ := \$v1975\(0 to 3);
                \$v1974\ := ""&\$v1975\(4);
                case \$v1976\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1972\ := \$arr1644_ptr_take\;
                if \$v1972\(0) = '1' then
                  state_var2247 <= q_wait1971;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1969;
                end if;
              when "0001" =>
                \$114_n\ := \$v1973\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1972\ := \$arr1644_ptr_take\;
                if \$v1972\(0) = '1' then
                  state_var2247 <= q_wait1971;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1969;
                end if;
              when "0000" =>
                \$115_b\ := \$v1973\(0 to 0);
                \$v1977\ := \$115_b\;
                if \$v1977\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1972\ := \$arr1644_ptr_take\;
                  if \$v1972\(0) = '1' then
                    state_var2247 <= q_wait1971;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1969;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1992 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v184\ := \$arr1644_value\;
              \$v1989\ := \$v184\;
              \$v1990\ := \$v1989\(0 to 3);
              \$v1984\ := \$v1989\(4 to 67);
              case \$v1990\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1983\ := \$arr1644_ptr_take\;
                if \$v1983\(0) = '1' then
                  state_var2247 <= q_wait1982;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1980;
                end if;
              when "0011" =>
                \$113_p\ := \$v1984\(0 to 4);
                \$v1986\ := \$113_p\;
                \$v1987\ := \$v1986\(0 to 3);
                \$v1985\ := ""&\$v1986\(4);
                case \$v1987\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1983\ := \$arr1644_ptr_take\;
                if \$v1983\(0) = '1' then
                  state_var2247 <= q_wait1982;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1980;
                end if;
              when "0001" =>
                \$114_n\ := \$v1984\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("stack["));
                
                eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v1983\ := \$arr1644_ptr_take\;
                if \$v1983\(0) = '1' then
                  state_var2247 <= q_wait1982;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                  state_var2247 <= pause_getI1980;
                end if;
              when "0000" =>
                \$115_b\ := \$v1984\(0 to 0);
                \$v1988\ := \$115_b\;
                if \$v1988\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1983\ := \$arr1644_ptr_take\;
                  if \$v1983\(0) = '1' then
                    state_var2247 <= q_wait1982;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                    state_var2247 <= pause_getI1980;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2000 =>
              \$arr1644_ptr_take\(0) := '0';
              \value\ := \$arr1644_value\;
              \$v1997\ := \value\;
              \$v1998\ := \$v1997\(0 to 3);
              \$v1743\ := \$v1997\(4 to 67);
              case \$v1998\ is
              when "0100" =>
                \$v1114\ := \$v1743\(0 to 63);
                \$v1756\ := \$arr1643_ptr_take\;
                if \$v1756\(0) = '1' then
                  state_var2247 <= q_wait1755;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$v1752\ := \$v1114\(32 to 63);
                  \$arr1643_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(32 to 63)));
                  \$arr1643_write_request\ <= '1';
                  \$arr1643_write\ <= "0001" & \$v1752\&X"00000000";
                  state_var2247 <= pause_setI1753;
                end if;
              when "0011" =>
                p := \$v1743\(0 to 4);
                \$v1995\ := p;
                \$v1996\ := \$v1995\(0 to 3);
                \$v1757\ := ""&\$v1995\(4);
                case \$v1996\ is
                when "0101" =>
                  \$v1782\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v1782\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2247 <= \$120_forever5481625\;
                  else
                    \$v1781\ := \$arr1644_ptr_take\;
                    if \$v1781\(0) = '1' then
                      state_var2247 <= q_wait1780;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                      state_var2247 <= pause_getI1778;
                    end if;
                  end if;
                when "0110" =>
                  \$v1843\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v1843\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2247 <= \$120_forever5481628\;
                  else
                    \$v1842\ := \$arr1644_ptr_take\;
                    if \$v1842\(0) = '1' then
                      state_var2247 <= q_wait1841;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2247 <= pause_getI1839;
                    end if;
                  end if;
                when "0100" =>
                  \$v1862\ := eclat_neq(\$192_n\ & "00000000000000000000000000000010");
                  if \$v1862\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut exactement 2 arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2247 <= \$120_forever5481631\;
                  else
                    \$v1861\ := \$arr1644_ptr_take\;
                    if \$v1861\(0) = '1' then
                      state_var2247 <= q_wait1860;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                      state_var2247 <= pause_getI1858;
                    end if;
                  end if;
                when "0011" =>
                  \$v1874\ := eclat_lt(\$192_n\ & "00000000000000000000000000000001");
                  if \$v1874\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("pas assez d'arguments"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2247 <= \$120_forever5481633\;
                  else
                    \$v1873\ := \$arr1644_ptr_take\;
                    if \$v1873\(0) = '1' then
                      state_var2247 <= q_wait1872;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                      state_var2247 <= pause_getI1870;
                    end if;
                  end if;
                when "0010" =>
                  \$146_mul544_arg\ := \$192_n\ & "00000000000000000000000000000001" & \$149_vm_run_code521_arg\(0 to 31);
                  state_var2247 <= \$146_mul544\;
                when "0001" =>
                  \$v1957\ := eclat_lt(\$192_n\ & "00000000000000000000000000000010");
                  if \$v1957\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("il faut 2 arguments pour la soustraction"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var2247 <= \$120_forever5481635\;
                  else
                    \$v1956\ := \$arr1644_ptr_take\;
                    if \$v1956\(0) = '1' then
                      state_var2247 <= q_wait1955;
                    else
                      \$arr1644_ptr_take\(0) := '1';
                      \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                      state_var2247 <= pause_getI1953;
                    end if;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("stack["));
                  
                  eclat_print_int(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001"));
                  
                  eclat_print_string(of_string("] <-"));
                  
                  \$v1994\ := \$arr1644_ptr_take\;
                  if \$v1994\(0) = '1' then
                    state_var2247 <= q_wait1993;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI1991;
                  end if;
                when others =>
                  \$165\ := \$149_vm_run_code521_arg\(0 to 293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                end case;
              when others =>
                \$165\ := \$149_vm_run_code521_arg\(0 to 293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              end case;
            when pause_getII2013 =>
              \$arr1647_ptr_take\(0) := '0';
              \$v1499\ := \$arr1647_value\;
              \$v2011\ := \$arr1644_ptr_take\;
              if \$v2011\(0) = '1' then
                state_var2247 <= q_wait2010;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$v1499\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= v;
                state_var2247 <= pause_setI2008;
              end if;
            when pause_getII2017 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2015\ := \$arr1647_ptr_take\;
              if \$v2015\(0) = '1' then
                state_var2247 <= q_wait2014;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(96 to 127)));
                state_var2247 <= pause_getI2012;
              end if;
            when pause_getII2024 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2021\ := v;
              \$v2022\ := \$v2021\(0 to 3);
              \$v2020\ := \$v2021\(4 to 67);
              case \$v2022\ is
              when "0000" =>
                x := \$v2020\(0 to 0);
                condition := x;
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & 
                eclat_if(condition & \$149_vm_run_code521_arg\(64 to 95) & eclat_sub(\$195_l\ & "00000000000000000000000000000001")) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when others =>
                condition := eclat_false;
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & 
                eclat_if(condition & \$149_vm_run_code521_arg\(64 to 95) & eclat_sub(\$195_l\ & "00000000000000000000000000000001")) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              end case;
            when pause_getII2031 =>
              \$arr1644_ptr_take\(0) := '0';
              v := \$arr1644_value\;
              \$v2028\ := v;
              \$v2029\ := \$v2028\(0 to 3);
              \$v2027\ := \$v2028\(4 to 67);
              case \$v2029\ is
              when "0000" =>
                x := \$v2027\(0 to 0);
                cond := x;
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$196_l\ & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(64 to 95)) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when others =>
                cond := eclat_false;
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & 
                eclat_if(cond & eclat_sub(\$196_l\ & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(64 to 95)) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              end case;
            when pause_getII2039 =>
              \$arr1644_ptr_take\(0) := '0';
              var := \$arr1644_value\;
              \$v2037\ := \$arr1643_ptr_take\;
              if \$v2037\(0) = '1' then
                state_var2247 <= q_wait2036;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$197_i\)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= var;
                state_var2247 <= pause_setI2034;
              end if;
            when pause_getII2047 =>
              \$arr1643_ptr_take\(0) := '0';
              local_value := \$arr1643_value\;
              \$v2045\ := \$arr1644_ptr_take\;
              if \$v2045\(0) = '1' then
                state_var2247 <= q_wait2044;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= local_value;
                state_var2247 <= pause_setI2042;
              end if;
            when pause_getII2058 =>
              \$arr1643_ptr_take\(0) := '0';
              \$v221\ := \$arr1643_value\;
              \$v2055\ := \$v221\;
              \$v2056\ := \$v2055\(0 to 3);
              \$v2050\ := \$v2055\(4 to 67);
              case \$v2056\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2247 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                  state_var2247 <= pause_getI2046;
                end if;
              when "0011" =>
                \$113_p\ := \$v2050\(0 to 4);
                \$v2052\ := \$113_p\;
                \$v2053\ := \$v2052\(0 to 3);
                \$v2051\ := ""&\$v2052\(4);
                case \$v2053\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2247 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                  state_var2247 <= pause_getI2046;
                end if;
              when "0001" =>
                \$114_n\ := \$v2050\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$v2049\ := \$arr1643_ptr_take\;
                if \$v2049\(0) = '1' then
                  state_var2247 <= q_wait2048;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                  state_var2247 <= pause_getI2046;
                end if;
              when "0000" =>
                \$115_b\ := \$v2050\(0 to 0);
                \$v2054\ := \$115_b\;
                if \$v2054\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$v2049\ := \$arr1643_ptr_take\;
                  if \$v2049\(0) = '1' then
                    state_var2247 <= q_wait2048;
                  else
                    \$arr1643_ptr_take\(0) := '1';
                    \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                    state_var2247 <= pause_getI2046;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2066 =>
              \$arr1645_ptr_take\(0) := '0';
              \$v225\ := \$arr1645_value\;
              \$v2064\ := \$arr1644_ptr_take\;
              if \$v2064\(0) = '1' then
                state_var2247 <= q_wait2063;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$v225\;
                state_var2247 <= pause_setI2061;
              end if;
            when pause_getII2074 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v229\ := \$arr1644_value\;
              \$v2072\ := \$arr1645_ptr_take\;
              if \$v2072\(0) = '1' then
                state_var2247 <= q_wait2071;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr_write\ <= to_integer(unsigned(\$201_i\));
                \$arr1645_write_request\ <= '1';
                \$arr1645_write\ <= \$v229\;
                state_var2247 <= pause_setI2069;
              end if;
            when pause_getII2085 =>
              \$arr1644_ptr_take\(0) := '0';
              \$v237\ := \$arr1644_value\;
              \$v2082\ := \$v237\;
              \$v2083\ := \$v2082\(0 to 3);
              \$v2077\ := \$v2082\(4 to 67);
              case \$v2083\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0011" =>
                \$113_p\ := \$v2077\(0 to 4);
                \$v2079\ := \$113_p\;
                \$v2080\ := \$v2079\(0 to 3);
                \$v2078\ := ""&\$v2079\(4);
                case \$v2080\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0001" =>
                \$114_n\ := \$v2077\(0 to 31);
                eclat_print_int(\$114_n\);
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0000" =>
                \$115_b\ := \$v2077\(0 to 0);
                \$v2081\ := \$115_b\;
                if \$v2081\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & eclat_true;
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII2096 =>
              \$arr1646_ptr_take\(0) := '0';
              \$191_instr\ := \$arr1646_value\;
              \$v2093\ := \$191_instr\;
              \$v2094\ := \$v2093\(0 to 3);
              \$v1742\ := \$v2093\(4 to 71);
              case \$v2094\ is
              when "1000" =>
                \$192_n\ := \$v1742\(0 to 31);
                \$v2002\ := \$arr1644_ptr_take\;
                if \$v2002\(0) = '1' then
                  state_var2247 <= q_wait2001;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI1999;
                end if;
              when "0110" =>
                \$193_l\ := \$v1742\(0 to 31);
                \$v2007\ := \$arr1644_ptr_take\;
                if \$v2007\(0) = '1' then
                  state_var2247 <= q_wait2006;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$v2003\ := \$193_l\ & \$149_vm_run_code521_arg\(32 to 63);
                  \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= "0100" & \$v2003\;
                  state_var2247 <= pause_setI2004;
                end if;
              when "1001" =>
                \$v2019\ := \$arr1644_ptr_take\;
                if \$v2019\(0) = '1' then
                  state_var2247 <= q_wait2018;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI2016;
                end if;
              when "1100" =>
                \$195_l\ := \$v1742\(0 to 31);
                \$v2026\ := \$arr1644_ptr_take\;
                if \$v2026\(0) = '1' then
                  state_var2247 <= q_wait2025;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI2023;
                end if;
              when "1011" =>
                \$196_l\ := \$v1742\(0 to 31);
                \$v2033\ := \$arr1644_ptr_take\;
                if \$v2033\(0) = '1' then
                  state_var2247 <= q_wait2032;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI2030;
                end if;
              when "0011" =>
                \$197_i\ := \$v1742\(0 to 31);
                \$v2041\ := \$arr1644_ptr_take\;
                if \$v2041\(0) = '1' then
                  state_var2247 <= q_wait2040;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI2038;
                end if;
              when "1010" =>
                \$198_l\ := \$v1742\(0 to 31);
                \$165\ := \$149_vm_run_code521_arg\(0 to 31) & \$149_vm_run_code521_arg\(32 to 63) & eclat_sub(\$198_l\ & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0100" =>
                \$199_i\ := \$v1742\(0 to 31);
                eclat_print_string(of_string("env "));
                
                eclat_print_int(\$149_vm_run_code521_arg\(32 to 63));
                
                eclat_print_newline(eclat_unit);
                
                eclat_print_string(of_string("Fetch["));
                
                eclat_print_int(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\));
                
                eclat_print_string(of_string("] <-"));
                
                \$v2060\ := \$arr1643_ptr_take\;
                if \$v2060\(0) = '1' then
                  state_var2247 <= q_wait2059;
                else
                  \$arr1643_ptr_take\(0) := '1';
                  \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                  state_var2247 <= pause_getI2057;
                end if;
              when "0010" =>
                \$200_i\ := \$v1742\(0 to 31);
                \$v2068\ := \$arr1645_ptr_take\;
                if \$v2068\(0) = '1' then
                  state_var2247 <= q_wait2067;
                else
                  \$arr1645_ptr_take\(0) := '1';
                  \$arr1645_ptr\ <= to_integer(unsigned(\$200_i\));
                  state_var2247 <= pause_getI2065;
                end if;
              when "0001" =>
                \$201_i\ := \$v1742\(0 to 31);
                \$v2076\ := \$arr1644_ptr_take\;
                if \$v2076\(0) = '1' then
                  state_var2247 <= q_wait2075;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                  state_var2247 <= pause_getI2073;
                end if;
              when "0000" =>
                \$165\ := \$149_vm_run_code521_arg\(0 to 31) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & eclat_add(\$149_vm_run_code521_arg\(128 to 159) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0111" =>
                \$v2088\ := eclat_eq(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & "00000000000000000000000000000000");
                if \$v2088\(0) = '1' then
                  \$v2087\ := \$arr1644_ptr_take\;
                  if \$v2087\(0) = '1' then
                    state_var2247 <= q_wait2086;
                  else
                    \$arr1644_ptr_take\(0) := '1';
                    \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                    state_var2247 <= pause_getI2084;
                  end if;
                else
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                end if;
              when "0101" =>
                \$204_v\ := \$v1742\(0 to 67);
                \$v2092\ := \$arr1644_ptr_take\;
                if \$v2092\(0) = '1' then
                  state_var2247 <= q_wait2091;
                else
                  \$arr1644_ptr_take\(0) := '1';
                  \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                  \$arr1644_write_request\ <= '1';
                  \$arr1644_write\ <= \$204_v\;
                  state_var2247 <= pause_setI2089;
                end if;
              when others =>
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var2247 <= \$208_forever5471620\;
              end case;
            when pause_setI1698 =>
              \$arr1643_write_request\ <= '0';
              state_var2247 <= pause_setII1699;
            when pause_setI1744 =>
              \$arr1647_write_request\ <= '0';
              state_var2247 <= pause_setII1745;
            when pause_setI1748 =>
              \$arr1647_write_request\ <= '0';
              state_var2247 <= pause_setII1749;
            when pause_setI1753 =>
              \$arr1643_write_request\ <= '0';
              state_var2247 <= pause_setII1754;
            when pause_setI1758 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1759;
            when pause_setI1792 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1793;
            when pause_setI1844 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1845;
            when pause_setI1863 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1864;
            when pause_setI1875 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1876;
            when pause_setI1913 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1914;
            when pause_setI1958 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII1959;
            when pause_setI2004 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII2005;
            when pause_setI2008 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII2009;
            when pause_setI2034 =>
              \$arr1643_write_request\ <= '0';
              state_var2247 <= pause_setII2035;
            when pause_setI2042 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII2043;
            when pause_setI2061 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII2062;
            when pause_setI2069 =>
              \$arr1645_write_request\ <= '0';
              state_var2247 <= pause_setII2070;
            when pause_setI2089 =>
              \$arr1644_write_request\ <= '0';
              state_var2247 <= pause_setII2090;
            when pause_setII1699 =>
              \$arr1643_ptr_take\(0) := '0';
              \$143_copy_args_to_heap518_arg\ := eclat_sub(\$143_copy_args_to_heap518_arg\(0 to 31) & "00000000000000000000000000000001") & \$143_copy_args_to_heap518_arg\(32 to 63) & eclat_add(\$143_copy_args_to_heap518_arg\(64 to 95) & "00000000000000000000000000000001");
              state_var2247 <= \$143_copy_args_to_heap518\;
            when pause_setII1745 =>
              \$arr1647_ptr_take\(0) := '0';
              \$165\ := eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(\$v1114\(32 to 63) & "00000000000000000000000000000001") & eclat_sub(\$v1114\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1749 =>
              \$arr1647_ptr_take\(0) := '0';
              \$v1747\ := \$arr1647_ptr_take\;
              if \$v1747\(0) = '1' then
                state_var2247 <= q_wait1746;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$v1114\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(96 to 127);
                state_var2247 <= pause_setI1744;
              end if;
            when pause_setII1754 =>
              \$arr1643_ptr_take\(0) := '0';
              \$143_copy_args_to_heap518_arg\ := \$192_n\ & \$149_vm_run_code521_arg\(0 to 31) & eclat_add(\$149_vm_run_code521_arg\(32 to 63) & "00000000000000000000000000000001");
              state_var2247 <= \$143_copy_args_to_heap518\;
            when pause_setII1759 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1793 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_string(of_string("ICIIIIIIIII"));
              
              \$v1790\ := eclat_gt(fst_operand & scd_operand);
              \$v1788\ := "0000" & \$v1790\&"000"& X"000000000000000";
              \$v1789\ := \$v1788\(0 to 3);
              \$v1783\ := \$v1788\(4 to 67);
              case \$v1789\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0011" =>
                \$113_p\ := \$v1783\(0 to 4);
                \$v1785\ := \$113_p\;
                \$v1786\ := \$v1785\(0 to 3);
                \$v1784\ := ""&\$v1785\(4);
                case \$v1786\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0001" =>
                \$114_n\ := \$v1783\(0 to 31);
                eclat_print_int(\$114_n\);
                
                eclat_print_newline(eclat_unit);
                
                \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                \$v1741\ := ""&\$165\(293);
                if \$v1741\(0) = '1' then
                  \$149_vm_run_code521_result\ := eclat_unit;
                  result1695 := \$149_vm_run_code521_result\;
                  rdy1696 := eclat_true;
                  state_var2247 <= compute1697;
                else
                  \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                  state_var2247 <= \$149_vm_run_code521\;
                end if;
              when "0000" =>
                \$115_b\ := \$v1783\(0 to 0);
                \$v1787\ := \$115_b\;
                if \$v1787\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
                  \$v1741\ := ""&\$165\(293);
                  if \$v1741\(0) = '1' then
                    \$149_vm_run_code521_result\ := eclat_unit;
                    result1695 := \$149_vm_run_code521_result\;
                    rdy1696 := eclat_true;
                    state_var2247 <= compute1697;
                  else
                    \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                    state_var2247 <= \$149_vm_run_code521\;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_setII1845 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1864 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1876 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1914 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_int(eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat));
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII1959 =>
              \$arr1644_ptr_take\(0) := '0';
              eclat_print_int(resultat);
              
              eclat_print_newline(eclat_unit);
              
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2005 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2009 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$v1499\(0 to 31) & "00000000000000000000000000000001") & \$v1499\(32 to 63) & \$v1499\(64 to 95) & \$v1499\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2035 =>
              \$arr1643_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2043 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2062 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2070 =>
              \$arr1645_ptr_take\(0) := '0';
              \$165\ := eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when pause_setII2090 =>
              \$arr1644_ptr_take\(0) := '0';
              \$165\ := eclat_add(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127) & \$149_vm_run_code521_arg\(128 to 159) & \$149_vm_run_code521_arg\(160 to 191) & \$149_vm_run_code521_arg\(192 to 292) & ""&\$149_vm_run_code521_arg\(293);
              \$v1741\ := ""&\$165\(293);
              if \$v1741\(0) = '1' then
                \$149_vm_run_code521_result\ := eclat_unit;
                result1695 := \$149_vm_run_code521_result\;
                rdy1696 := eclat_true;
                state_var2247 <= compute1697;
              else
                \$149_vm_run_code521_arg\ := \$165\(0 to 31) & \$165\(32 to 63) & eclat_add(\$165\(64 to 95) & "00000000000000000000000000000001") & \$165\(96 to 127) & \$165\(128 to 159) & \$165\(160 to 191) & \$165\(192 to 292) & ""&\$165\(293) & ""&\$149_vm_run_code521_arg\(294);
                state_var2247 <= \$149_vm_run_code521\;
              end if;
            when q_wait1700 =>
              \$v1701\ := \$arr1643_ptr_take\;
              if \$v1701\(0) = '1' then
                state_var2247 <= q_wait1700;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(\$143_copy_args_to_heap518_arg\(64 to 95)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= \$389\;
                state_var2247 <= pause_setI1698;
              end if;
            when q_wait1704 =>
              \$v1705\ := \$arr1644_ptr_take\;
              if \$v1705\(0) = '1' then
                state_var2247 <= q_wait1704;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$143_copy_args_to_heap518_arg\(32 to 63) & \$143_copy_args_to_heap518_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1702;
              end if;
            when q_wait1714 =>
              \$v1715\ := \$arr1644_ptr_take\;
              if \$v1715\(0) = '1' then
                state_var2247 <= q_wait1714;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$145_div543_arg\(64 to 95) & "00000000000000000000000000000001") & \$145_div543_arg\(0 to 31))));
                state_var2247 <= pause_getI1712;
              end if;
            when q_wait1722 =>
              \$v1723\ := \$arr1644_ptr_take\;
              if \$v1723\(0) = '1' then
                state_var2247 <= q_wait1722;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$146_mul544_arg\(64 to 95) & "00000000000000000000000000000001") & \$146_mul544_arg\(0 to 31))));
                state_var2247 <= pause_getI1720;
              end if;
            when q_wait1730 =>
              \$v1731\ := \$arr1644_ptr_take\;
              if \$v1731\(0) = '1' then
                state_var2247 <= q_wait1730;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$147_sub545_arg\(64 to 95) & "00000000000000000000000000000001") & \$147_sub545_arg\(0 to 31))));
                state_var2247 <= pause_getI1728;
              end if;
            when q_wait1738 =>
              \$v1739\ := \$arr1644_ptr_take\;
              if \$v1739\(0) = '1' then
                state_var2247 <= q_wait1738;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$148_add546_arg\(64 to 95) & "00000000000000000000000000000001") & \$148_add546_arg\(0 to 31))));
                state_var2247 <= pause_getI1736;
              end if;
            when q_wait1746 =>
              \$v1747\ := \$arr1647_ptr_take\;
              if \$v1747\(0) = '1' then
                state_var2247 <= q_wait1746;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(96 to 127) & "00000000000000000000000000000001")));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & eclat_add(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$192_n\) & "00000000000000000000000000000001") & eclat_sub(\$v1114\(0 to 31) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(96 to 127);
                state_var2247 <= pause_setI1744;
              end if;
            when q_wait1750 =>
              \$v1751\ := \$arr1647_ptr_take\;
              if \$v1751\(0) = '1' then
                state_var2247 <= q_wait1750;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(96 to 127)));
                \$arr1647_write_request\ <= '1';
                \$arr1647_write\ <= eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001") & \$149_vm_run_code521_arg\(32 to 63) & \$149_vm_run_code521_arg\(64 to 95) & \$149_vm_run_code521_arg\(96 to 127);
                state_var2247 <= pause_setI1748;
              end if;
            when q_wait1755 =>
              \$v1756\ := \$arr1643_ptr_take\;
              if \$v1756\(0) = '1' then
                state_var2247 <= q_wait1755;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$v1752\ := \$v1114\(32 to 63);
                \$arr1643_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(32 to 63)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= "0001" & \$v1752\&X"00000000";
                state_var2247 <= pause_setI1753;
              end if;
            when q_wait1760 =>
              \$v1761\ := \$arr1644_ptr_take\;
              if \$v1761\(0) = '1' then
                state_var2247 <= q_wait1760;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001") & \$192_n\)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0000" & res&"000"& X"000000000000000";
                state_var2247 <= pause_setI1758;
              end if;
            when q_wait1776 =>
              \$v1777\ := \$arr1644_ptr_take\;
              if \$v1777\(0) = '1' then
                state_var2247 <= q_wait1776;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2247 <= pause_getI1774;
              end if;
            when q_wait1780 =>
              \$v1781\ := \$arr1644_ptr_take\;
              if \$v1781\(0) = '1' then
                state_var2247 <= q_wait1780;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2247 <= pause_getI1778;
              end if;
            when q_wait1794 =>
              \$v1795\ := \$arr1644_ptr_take\;
              if \$v1795\(0) = '1' then
                state_var2247 <= q_wait1794;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v1791\ := eclat_gt(fst_operand & scd_operand);
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0000" & \$v1791\&"000"& X"000000000000000";
                state_var2247 <= pause_setI1792;
              end if;
            when q_wait1805 =>
              \$v1806\ := \$arr1644_ptr_take\;
              if \$v1806\(0) = '1' then
                state_var2247 <= q_wait1805;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1803;
              end if;
            when q_wait1816 =>
              \$v1817\ := \$arr1644_ptr_take\;
              if \$v1817\(0) = '1' then
                state_var2247 <= q_wait1816;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2247 <= pause_getI1814;
              end if;
            when q_wait1827 =>
              \$v1828\ := \$arr1644_ptr_take\;
              if \$v1828\(0) = '1' then
                state_var2247 <= q_wait1827;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2247 <= pause_getI1825;
              end if;
            when q_wait1834 =>
              \$v1835\ := \$arr1644_ptr_take\;
              if \$v1835\(0) = '1' then
                state_var2247 <= q_wait1834;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2247 <= pause_getI1832;
              end if;
            when q_wait1841 =>
              \$v1842\ := \$arr1644_ptr_take\;
              if \$v1842\(0) = '1' then
                state_var2247 <= q_wait1841;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2247 <= pause_getI1839;
              end if;
            when q_wait1846 =>
              \$v1847\ := \$arr1644_ptr_take\;
              if \$v1847\(0) = '1' then
                state_var2247 <= q_wait1846;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2247 <= pause_setI1844;
              end if;
            when q_wait1853 =>
              \$v1854\ := \$arr1644_ptr_take\;
              if \$v1854\(0) = '1' then
                state_var2247 <= q_wait1853;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000010")));
                state_var2247 <= pause_getI1851;
              end if;
            when q_wait1860 =>
              \$v1861\ := \$arr1644_ptr_take\;
              if \$v1861\(0) = '1' then
                state_var2247 <= q_wait1860;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000011")));
                state_var2247 <= pause_getI1858;
              end if;
            when q_wait1865 =>
              \$v1866\ := \$arr1644_ptr_take\;
              if \$v1866\(0) = '1' then
                state_var2247 <= q_wait1865;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2247 <= pause_setI1863;
              end if;
            when q_wait1872 =>
              \$v1873\ := \$arr1644_ptr_take\;
              if \$v1873\(0) = '1' then
                state_var2247 <= q_wait1872;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1870;
              end if;
            when q_wait1877 =>
              \$v1878\ := \$arr1644_ptr_take\;
              if \$v1878\(0) = '1' then
                state_var2247 <= q_wait1877;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2247 <= pause_setI1875;
              end if;
            when q_wait1888 =>
              \$v1889\ := \$arr1644_ptr_take\;
              if \$v1889\(0) = '1' then
                state_var2247 <= q_wait1888;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1886;
              end if;
            when q_wait1899 =>
              \$v1900\ := \$arr1644_ptr_take\;
              if \$v1900\(0) = '1' then
                state_var2247 <= q_wait1899;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                state_var2247 <= pause_getI1897;
              end if;
            when q_wait1910 =>
              \$v1911\ := \$arr1644_ptr_take\;
              if \$v1911\(0) = '1' then
                state_var2247 <= q_wait1910;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1908;
              end if;
            when q_wait1915 =>
              \$v1916\ := \$arr1644_ptr_take\;
              if \$v1916\(0) = '1' then
                state_var2247 <= q_wait1915;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v1912\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & \$v1912\&X"00000000";
                state_var2247 <= pause_setI1913;
              end if;
            when q_wait1926 =>
              \$v1927\ := \$arr1644_ptr_take\;
              if \$v1927\(0) = '1' then
                state_var2247 <= q_wait1926;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1924;
              end if;
            when q_wait1937 =>
              \$v1938\ := \$arr1644_ptr_take\;
              if \$v1938\(0) = '1' then
                state_var2247 <= q_wait1937;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                state_var2247 <= pause_getI1935;
              end if;
            when q_wait1948 =>
              \$v1949\ := \$arr1644_ptr_take\;
              if \$v1949\(0) = '1' then
                state_var2247 <= q_wait1948;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1946;
              end if;
            when q_wait1955 =>
              \$v1956\ := \$arr1644_ptr_take\;
              if \$v1956\(0) = '1' then
                state_var2247 <= q_wait1955;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1953;
              end if;
            when q_wait1960 =>
              \$v1961\ := \$arr1644_ptr_take\;
              if \$v1961\(0) = '1' then
                state_var2247 <= q_wait1960;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0001" & resultat&X"00000000";
                state_var2247 <= pause_setI1958;
              end if;
            when q_wait1971 =>
              \$v1972\ := \$arr1644_ptr_take\;
              if \$v1972\(0) = '1' then
                state_var2247 <= q_wait1971;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_add(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1969;
              end if;
            when q_wait1982 =>
              \$v1983\ := \$arr1644_ptr_take\;
              if \$v1983\(0) = '1' then
                state_var2247 <= q_wait1982;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\)));
                state_var2247 <= pause_getI1980;
              end if;
            when q_wait1993 =>
              \$v1994\ := \$arr1644_ptr_take\;
              if \$v1994\(0) = '1' then
                state_var2247 <= q_wait1993;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & \$192_n\) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1991;
              end if;
            when q_wait2001 =>
              \$v2002\ := \$arr1644_ptr_take\;
              if \$v2002\(0) = '1' then
                state_var2247 <= q_wait2001;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI1999;
              end if;
            when q_wait2006 =>
              \$v2007\ := \$arr1644_ptr_take\;
              if \$v2007\(0) = '1' then
                state_var2247 <= q_wait2006;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$v2003\ := \$193_l\ & \$149_vm_run_code521_arg\(32 to 63);
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= "0100" & \$v2003\;
                state_var2247 <= pause_setI2004;
              end if;
            when q_wait2010 =>
              \$v2011\ := \$arr1644_ptr_take\;
              if \$v2011\(0) = '1' then
                state_var2247 <= q_wait2010;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$v1499\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= v;
                state_var2247 <= pause_setI2008;
              end if;
            when q_wait2014 =>
              \$v2015\ := \$arr1647_ptr_take\;
              if \$v2015\(0) = '1' then
                state_var2247 <= q_wait2014;
              else
                \$arr1647_ptr_take\(0) := '1';
                \$arr1647_ptr\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(96 to 127)));
                state_var2247 <= pause_getI2012;
              end if;
            when q_wait2018 =>
              \$v2019\ := \$arr1644_ptr_take\;
              if \$v2019\(0) = '1' then
                state_var2247 <= q_wait2018;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2016;
              end if;
            when q_wait2025 =>
              \$v2026\ := \$arr1644_ptr_take\;
              if \$v2026\(0) = '1' then
                state_var2247 <= q_wait2025;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2023;
              end if;
            when q_wait2032 =>
              \$v2033\ := \$arr1644_ptr_take\;
              if \$v2033\(0) = '1' then
                state_var2247 <= q_wait2032;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2030;
              end if;
            when q_wait2036 =>
              \$v2037\ := \$arr1643_ptr_take\;
              if \$v2037\(0) = '1' then
                state_var2247 <= q_wait2036;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr_write\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$197_i\)));
                \$arr1643_write_request\ <= '1';
                \$arr1643_write\ <= var;
                state_var2247 <= pause_setI2034;
              end if;
            when q_wait2040 =>
              \$v2041\ := \$arr1644_ptr_take\;
              if \$v2041\(0) = '1' then
                state_var2247 <= q_wait2040;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2038;
              end if;
            when q_wait2044 =>
              \$v2045\ := \$arr1644_ptr_take\;
              if \$v2045\(0) = '1' then
                state_var2247 <= q_wait2044;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= local_value;
                state_var2247 <= pause_setI2042;
              end if;
            when q_wait2048 =>
              \$v2049\ := \$arr1643_ptr_take\;
              if \$v2049\(0) = '1' then
                state_var2247 <= q_wait2048;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                state_var2247 <= pause_getI2046;
              end if;
            when q_wait2059 =>
              \$v2060\ := \$arr1643_ptr_take\;
              if \$v2060\(0) = '1' then
                state_var2247 <= q_wait2059;
              else
                \$arr1643_ptr_take\(0) := '1';
                \$arr1643_ptr\ <= to_integer(unsigned(eclat_add(\$149_vm_run_code521_arg\(32 to 63) & \$199_i\)));
                state_var2247 <= pause_getI2057;
              end if;
            when q_wait2063 =>
              \$v2064\ := \$arr1644_ptr_take\;
              if \$v2064\(0) = '1' then
                state_var2247 <= q_wait2063;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$v225\;
                state_var2247 <= pause_setI2061;
              end if;
            when q_wait2067 =>
              \$v2068\ := \$arr1645_ptr_take\;
              if \$v2068\(0) = '1' then
                state_var2247 <= q_wait2067;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr\ <= to_integer(unsigned(\$200_i\));
                state_var2247 <= pause_getI2065;
              end if;
            when q_wait2071 =>
              \$v2072\ := \$arr1645_ptr_take\;
              if \$v2072\(0) = '1' then
                state_var2247 <= q_wait2071;
              else
                \$arr1645_ptr_take\(0) := '1';
                \$arr1645_ptr_write\ <= to_integer(unsigned(\$201_i\));
                \$arr1645_write_request\ <= '1';
                \$arr1645_write\ <= \$v229\;
                state_var2247 <= pause_setI2069;
              end if;
            when q_wait2075 =>
              \$v2076\ := \$arr1644_ptr_take\;
              if \$v2076\(0) = '1' then
                state_var2247 <= q_wait2075;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2073;
              end if;
            when q_wait2086 =>
              \$v2087\ := \$arr1644_ptr_take\;
              if \$v2087\(0) = '1' then
                state_var2247 <= q_wait2086;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr\ <= to_integer(unsigned(eclat_sub(\$149_vm_run_code521_arg\(0 to 31) & "00000000000000000000000000000001")));
                state_var2247 <= pause_getI2084;
              end if;
            when q_wait2091 =>
              \$v2092\ := \$arr1644_ptr_take\;
              if \$v2092\(0) = '1' then
                state_var2247 <= q_wait2091;
              else
                \$arr1644_ptr_take\(0) := '1';
                \$arr1644_ptr_write\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(0 to 31)));
                \$arr1644_write_request\ <= '1';
                \$arr1644_write\ <= \$204_v\;
                state_var2247 <= pause_setI2089;
              end if;
            when q_wait2097 =>
              \$v2098\ := \$arr1646_ptr_take\;
              if \$v2098\(0) = '1' then
                state_var2247 <= q_wait2097;
              else
                \$arr1646_ptr_take\(0) := '1';
                \$arr1646_ptr\ <= to_integer(unsigned(\$149_vm_run_code521_arg\(64 to 95)));
                state_var2247 <= pause_getI2095;
              end if;
            when compute1697 =>
              rdy1696 := eclat_false;
              eclat_print_string(of_string("START (cy="));
              
              eclat_print_int(\$135_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              \$v2100\ := eclat_unit;
              \$149_vm_run_code521_arg\ := "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & eclat_false & "00000000000000000000000000000000" & "0010" & \$v2100\&"000"& X"000000000000000" & eclat_false & argument;
              state_var2247 <= \$149_vm_run_code521\;
            end case;
            \$v2102\ := eclat_not(rdy1696);
            if \$v2102\(0) = '1' then
              result1695 := eclat_unit;
            end if;
            \$136\ := result1695 & rdy1696;
            \$v1694\ := ""&\$136\(1);
            if \$v1694\(0) = '1' then
              eclat_print_string(of_string("END (cy="));
              
              eclat_print_int(\$135_cy\);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              result1648 := eclat_unit;
              eclat_print_newline(eclat_unit);
              
              rdy1649 := eclat_true;
              \state\ <= compute1650;
            else
              result1648 := eclat_unit;
              rdy1649 := eclat_true;
              \state\ <= compute1650;
            end if;
          end case;
          
          result <= result1648;
          rdy <= rdy1649;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
